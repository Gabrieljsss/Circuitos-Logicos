CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 181 342 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21488 90
2 5V
6 4 20 12
2 B5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
364 0 0
2
5.89819e-315 5.34643e-315
0
13 Logic Switch~
5 214 342 0 1 11
0 34
0
0 0 21360 90
2 0V
10 0 24 8
2 B4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3656 0 0
2
5.89819e-315 5.32571e-315
0
13 Logic Switch~
5 246 342 0 1 11
0 33
0
0 0 21488 90
2 0V
11 0 25 8
2 B3
9 -9 23 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3131 0 0
2
5.89819e-315 5.30499e-315
0
13 Logic Switch~
5 277 342 0 1 11
0 32
0
0 0 21488 90
2 0V
9 -1 23 7
2 B2
10 -11 24 -3
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6772 0 0
2
5.89819e-315 5.26354e-315
0
13 Logic Switch~
5 96 347 0 1 11
0 5
0
0 0 21360 90
2 0V
11 0 25 8
2 B1
7 -9 21 -1
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9557 0 0
2
5.89819e-315 0
0
13 Logic Switch~
5 59 91 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 A1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5789 0 0
2
5.89819e-315 0
0
13 Logic Switch~
5 192 90 0 1 11
0 38
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 A5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7328 0 0
2
5.89819e-315 0
0
13 Logic Switch~
5 211 91 0 1 11
0 37
0
0 0 21360 270
2 0V
-6 -22 8 -14
2 A4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4799 0 0
2
5.89819e-315 0
0
13 Logic Switch~
5 231 91 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-8 -21 6 -13
2 A3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9196 0 0
2
5.89819e-315 0
0
13 Logic Switch~
5 249 91 0 1 11
0 39
0
0 0 21488 270
2 0V
-5 -20 9 -12
2 A2
-7 -31 7 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3857 0 0
2
5.89819e-315 0
0
6 74136~
219 472 372 0 3 22
0 7 5 3
0
0 0 624 0
7 74LS136
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7125 0 0
2
43023.6 0
0
9 2-In AND~
219 553 317 0 3 22
0 3 4 6
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3641 0 0
2
43023.6 0
0
9 Inverter~
13 490 230 0 2 22
0 7 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
9821 0 0
2
43023.6 0
0
7 Ground~
168 746 107 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3187 0 0
2
43023.5 0
0
9 CC 7-Seg~
183 1019 97 0 17 19
10 17 18 19 20 21 22 23 44 2
1 1 1 1 1 1 0 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
762 0 0
2
43023.5 0
0
9 CC 7-Seg~
183 1119 98 0 17 19
10 25 26 27 28 29 30 31 45 2
0 1 1 0 0 1 1 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
39 0 0
2
5.89819e-315 0
0
6 74LS48
188 917 203 0 14 29
0 12 11 10 9 46 47 31 30 29
28 27 26 25 48
0
0 0 4336 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9450 0 0
2
5.89819e-315 0
0
6 74LS48
188 918 326 0 14 29
0 2 2 2 6 49 50 23 22 21
20 19 18 17 51
0
0 0 4336 0
7 74LS248
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3236 0 0
2
5.89819e-315 0
0
6 74LS83
105 809 176 0 14 29
0 8 2 8 2 16 15 14 13 2
12 11 10 9 52
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U4
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3321 0 0
2
5.89819e-315 0
0
2 +V
167 337 271 0 1 3
0 24
0
0 0 53488 180
2 5V
9 -2 23 6
2 V1
8 -12 22 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8879 0 0
2
5.89819e-315 0
0
7 Ground~
168 1067 33 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5433 0 0
2
5.89819e-315 0
0
9 Inverter~
13 275 281 0 2 22
0 32 43
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U3D
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
3679 0 0
2
5.89819e-315 0
0
9 Inverter~
13 244 281 0 2 22
0 33 42
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U3C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
9342 0 0
2
5.89819e-315 0
0
9 Inverter~
13 212 281 0 2 22
0 34 41
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U3B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3623 0 0
2
5.89819e-315 0
0
9 Inverter~
13 179 281 0 2 22
0 35 40
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U3A
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3722 0 0
2
5.89819e-315 0
0
6 74LS83
105 397 185 0 14 29
0 38 37 36 39 40 41 42 43 24
16 15 14 13 7
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U2
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
8993 0 0
2
5.89819e-315 5.26354e-315
0
51
3 1 3 0 0 4224 0 11 12 0 0 3
505 372
505 308
529 308
2 1 4 0 0 8320 0 12 6 0 0 4
529 326
529 465
59 465
59 103
1 2 5 0 0 8320 0 5 11 0 0 5
97 334
97 311
420 311
420 381
456 381
3 4 6 0 0 4224 0 12 18 0 0 2
574 317
886 317
0 1 7 0 0 4224 0 0 11 14 0 3
446 230
446 363
456 363
3 0 8 0 0 4096 0 19 0 0 7 2
777 158
715 158
2 1 8 0 0 4224 0 13 19 0 0 4
511 230
715 230
715 140
777 140
2 0 2 0 0 4096 0 19 0 0 13 2
777 149
746 149
1 0 2 0 0 4224 0 18 0 0 11 2
886 290
746 290
2 0 2 0 0 0 0 18 0 0 11 2
886 299
746 299
3 0 2 0 0 0 0 18 0 0 13 3
886 308
746 308
746 221
4 0 2 0 0 0 0 19 0 0 13 2
777 167
746 167
1 9 2 0 0 0 0 14 19 0 0 3
746 115
746 221
777 221
14 1 7 0 0 128 0 26 13 0 0 2
429 230
475 230
4 13 9 0 0 4224 0 17 19 0 0 2
885 194
841 194
3 12 10 0 0 4224 0 17 19 0 0 2
885 185
841 185
2 11 11 0 0 4224 0 17 19 0 0 2
885 176
841 176
1 10 12 0 0 4224 0 17 19 0 0 2
885 167
841 167
8 13 13 0 0 4224 0 19 26 0 0 2
777 203
429 203
7 12 14 0 0 4224 0 19 26 0 0 2
777 194
429 194
6 11 15 0 0 4224 0 19 26 0 0 2
777 185
429 185
5 10 16 0 0 4224 0 19 26 0 0 2
777 176
429 176
13 1 17 0 0 8320 0 18 15 0 0 3
950 344
998 344
998 133
2 12 18 0 0 4224 0 15 18 0 0 3
1004 133
1004 335
950 335
3 11 19 0 0 4224 0 15 18 0 0 3
1010 133
1010 326
950 326
4 10 20 0 0 4224 0 15 18 0 0 3
1016 133
1016 317
950 317
5 9 21 0 0 4224 0 15 18 0 0 3
1022 133
1022 308
950 308
8 6 22 0 0 8320 0 18 15 0 0 3
950 299
1028 299
1028 133
7 7 23 0 0 8320 0 18 15 0 0 3
950 290
1034 290
1034 133
9 1 2 0 0 0 0 15 21 0 0 3
1019 55
1019 41
1067 41
1 9 2 0 0 128 0 21 16 0 0 3
1067 41
1119 41
1119 56
9 1 24 0 0 4224 0 26 20 0 0 3
365 230
337 230
337 256
1 13 25 0 0 8320 0 16 17 0 0 3
1098 134
1098 221
949 221
2 12 26 0 0 8320 0 16 17 0 0 3
1104 134
1104 212
949 212
3 11 27 0 0 8320 0 16 17 0 0 3
1110 134
1110 203
949 203
10 4 28 0 0 4224 0 17 16 0 0 3
949 194
1116 194
1116 134
9 5 29 0 0 4224 0 17 16 0 0 3
949 185
1122 185
1122 134
8 6 30 0 0 4224 0 17 16 0 0 3
949 176
1128 176
1128 134
7 7 31 0 0 4224 0 17 16 0 0 3
949 167
1134 167
1134 134
1 1 32 0 0 4224 0 22 4 0 0 2
278 299
278 329
1 1 33 0 0 4224 0 23 3 0 0 2
247 299
247 329
1 1 34 0 0 4224 0 24 2 0 0 2
215 299
215 329
1 1 35 0 0 4224 0 25 1 0 0 2
182 299
182 329
3 1 36 0 0 4224 0 26 9 0 0 3
365 167
231 167
231 103
2 1 37 0 0 4224 0 26 8 0 0 3
365 158
211 158
211 103
1 1 38 0 0 8320 0 7 26 0 0 3
192 102
192 149
365 149
4 1 39 0 0 4224 0 26 10 0 0 3
365 176
249 176
249 103
5 2 40 0 0 4224 0 26 25 0 0 3
365 185
182 185
182 263
6 2 41 0 0 4224 0 26 24 0 0 3
365 194
215 194
215 263
7 2 42 0 0 4224 0 26 23 0 0 3
365 203
247 203
247 263
8 2 43 0 0 4224 0 26 22 0 0 3
365 212
278 212
278 263
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
197 364 288 385
206 371 278 386
9 2� D�gito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
66 364 155 385
74 371 146 386
9 1� D�gito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
18 35 107 56
26 42 98 57
9 1� D�gito
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
176 35 267 56
185 42 257 57
9 2� D�gito
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
