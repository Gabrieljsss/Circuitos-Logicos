CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1120 30 110 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
57
9 Inverter~
13 308 1780 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U11B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
6691 0 0
2
43361.4 0
0
9 Inverter~
13 310 1711 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U11A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
3551 0 0
2
43361.4 0
0
9 Inverter~
13 319 1648 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
3706 0 0
2
43361.4 0
0
9 Inverter~
13 321 1606 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
3136 0 0
2
43361.4 0
0
14 Logic Display~
6 680 1618 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3128 0 0
2
43361.4 0
0
8 4-In OR~
219 649 1635 0 1 22
0 0
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
5719 0 0
2
43361.4 0
0
5 4081~
219 420 1619 0 3 22
0 9 8 7
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
3268 0 0
2
43361.4 0
0
5 4081~
219 420 1543 0 3 22
0 9 8 7
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
9751 0 0
2
43361.4 0
0
9 Inverter~
13 285 1522 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
8844 0 0
2
43361.4 0
0
13 Logic Switch~
5 134 1711 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3948 0 0
2
43361.4 1
0
13 Logic Switch~
5 136 1788 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6695 0 0
2
43361.4 0
0
13 Logic Switch~
5 136 1662 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
429 0 0
2
43361.4 2
0
13 Logic Switch~
5 134 1585 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9630 0 0
2
43361.4 1
0
13 Logic Switch~
5 136 1521 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5453 0 0
2
43361.4 0
0
13 Logic Switch~
5 427 1980 0 1 11
0 6
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3703 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 429 1916 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8886 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 135 1221 0 1 11
0 9
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3762 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 133 1285 0 1 11
0 10
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
320 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 135 1362 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9974 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 121 938 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4655 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 119 861 0 1 11
0 17
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4985 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 121 797 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6515 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 120 626 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8791 0 0
2
43361.4 0
0
13 Logic Switch~
5 119 417 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
345 0 0
2
43361.4 1
0
13 Logic Switch~
5 117 481 0 1 11
0 34
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
43361.4 2
0
13 Logic Switch~
5 119 558 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8900 0 0
2
43361.4 3
0
13 Logic Switch~
5 119 281 0 1 11
0 36
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8368 0 0
2
43361.4 4
0
13 Logic Switch~
5 117 204 0 1 11
0 37
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3392 0 0
2
43361.4 5
0
13 Logic Switch~
5 119 140 0 1 11
0 39
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
851 0 0
2
43361.4 6
0
14 Logic Display~
6 658 1954 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8736 0 0
2
5.89862e-315 0
0
5 4081~
219 638 1971 0 3 22
0 4 3 2
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
593 0 0
2
5.89862e-315 0
0
5 4071~
219 507 2028 0 3 22
0 5 6 3
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
5432 0 0
2
5.89862e-315 0
0
5 4011~
219 524 1940 0 3 22
0 5 6 4
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 8 0
1 U
3595 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 537 1211 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3394 0 0
2
5.89862e-315 0
0
9 Inverter~
13 289 1365 0 2 22
0 12 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
9850 0 0
2
5.89862e-315 0
0
5 4071~
219 394 1320 0 3 22
0 10 11 8
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
9350 0 0
2
5.89862e-315 0
0
5 4081~
219 517 1229 0 3 22
0 9 8 7
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
9109 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 709 839 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7363 0 0
2
5.89862e-315 0
0
9 Inverter~
13 460 1023 0 2 22
0 17 18
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
570 0 0
2
5.89862e-315 0
0
8 3-In OR~
219 677 855 0 4 22
0 16 15 14 13
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U4B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 4 0
1 U
3544 0 0
2
5.89862e-315 0
0
5 4081~
219 500 1014 0 3 22
0 19 18 14
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
4354 0 0
2
5.89862e-315 0
0
5 4081~
219 495 870 0 3 22
0 17 20 15
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
563 0 0
2
5.89862e-315 0
0
5 4081~
219 499 751 0 3 22
0 22 21 16
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3846 0 0
2
5.89862e-315 0
0
9 Inverter~
13 290 933 0 2 22
0 20 21
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
3884 0 0
2
5.89862e-315 0
0
9 Inverter~
13 279 793 0 2 22
0 19 22
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
6770 0 0
2
5.89862e-315 0
0
14 Logic Display~
6 677 470 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6353 0 0
2
5.89862e-315 0
0
8 3-In OR~
219 645 487 0 4 22
0 26 25 24 23
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
8785 0 0
2
5.89862e-315 0
0
9 Inverter~
13 327 348 0 2 22
0 30 29
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3868 0 0
2
43361.4 7
0
9 3-In AND~
219 433 354 0 4 22
0 29 28 27 26
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 3 0
1 U
3562 0 0
2
43361.4 8
0
9 3-In AND~
219 439 449 0 4 22
0 30 28 31 25
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 1 0
1 U
3338 0 0
2
43361.4 9
0
9 3-In AND~
219 440 593 0 4 22
0 28 32 31 24
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 1 0
1 U
9932 0 0
2
43361.4 10
0
9 Inverter~
13 320 620 0 2 22
0 27 31
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
387 0 0
2
43361.4 11
0
9 Inverter~
13 315 542 0 2 22
0 33 32
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
5673 0 0
2
43361.4 12
0
9 Inverter~
13 320 471 0 2 22
0 34 28
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
4882 0 0
2
43361.4 13
0
14 Logic Display~
6 313 167 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3606 0 0
2
43361.4 14
0
9 Inverter~
13 193 145 0 2 22
0 39 38
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3577 0 0
2
43361.4 15
0
9 3-In AND~
219 292 184 0 4 22
0 38 37 36 35
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 1 0
1 U
6283 0 0
2
43361.4 16
0
64
2 4 0 0 0 0 0 1 6 0 0 4
329 1780
619 1780
619 1649
632 1649
1 1 0 0 0 0 0 11 1 0 0 4
148 1788
285 1788
285 1780
293 1780
2 3 0 0 0 0 0 2 6 0 0 4
331 1711
624 1711
624 1640
632 1640
1 1 0 0 0 0 0 10 2 0 0 2
146 1711
295 1711
3 2 0 0 0 0 0 7 6 0 0 4
441 1619
619 1619
619 1631
632 1631
3 1 0 0 0 0 0 8 6 0 0 4
441 1543
624 1543
624 1622
632 1622
2 2 0 0 0 0 0 3 7 0 0 4
340 1648
388 1648
388 1628
396 1628
1 1 0 0 0 0 0 12 3 0 0 3
148 1662
304 1662
304 1648
2 1 0 0 0 0 0 4 7 0 0 3
342 1606
396 1606
396 1610
0 1 0 0 0 0 0 0 4 11 0 3
260 1585
260 1606
306 1606
1 2 0 0 0 0 0 13 8 0 0 4
146 1585
388 1585
388 1552
396 1552
2 1 0 0 0 0 0 9 8 0 0 4
306 1522
388 1522
388 1534
396 1534
1 1 0 0 0 0 0 14 9 0 0 4
148 1521
262 1521
262 1522
270 1522
1 5 0 0 0 0 0 5 6 0 0 3
680 1636
680 1635
682 1635
1 3 2 0 0 4224 0 30 31 0 0 3
658 1972
658 1971
659 1971
2 3 3 0 0 4224 0 31 32 0 0 4
614 1980
548 1980
548 2028
540 2028
3 1 4 0 0 4224 0 33 31 0 0 4
551 1940
606 1940
606 1962
614 1962
0 1 5 0 0 4224 0 0 32 21 0 3
467 1916
467 2019
494 2019
0 2 6 0 0 4224 0 0 32 20 0 3
446 1980
446 2037
494 2037
1 2 6 0 0 0 0 15 33 0 0 4
439 1980
492 1980
492 1949
500 1949
1 1 5 0 0 0 0 16 33 0 0 3
441 1916
500 1916
500 1931
1 3 7 0 0 4224 0 34 37 0 0 2
537 1229
538 1229
3 2 8 0 0 8320 0 36 37 0 0 4
427 1320
485 1320
485 1238
493 1238
1 1 9 0 0 4224 0 17 37 0 0 4
147 1221
485 1221
485 1220
493 1220
1 1 10 0 0 4224 0 18 36 0 0 4
145 1285
373 1285
373 1311
381 1311
2 2 11 0 0 4224 0 35 36 0 0 4
310 1365
373 1365
373 1329
381 1329
1 1 12 0 0 4224 0 19 35 0 0 4
147 1362
266 1362
266 1365
274 1365
1 4 13 0 0 4224 0 38 40 0 0 3
709 857
709 855
710 855
3 3 14 0 0 8320 0 41 40 0 0 4
521 1014
651 1014
651 864
664 864
3 2 15 0 0 4224 0 42 40 0 0 4
516 870
656 870
656 855
665 855
3 1 16 0 0 4224 0 43 40 0 0 4
520 751
656 751
656 846
664 846
0 1 17 0 0 8192 0 0 39 37 0 3
164 861
164 1023
445 1023
2 2 18 0 0 4224 0 39 41 0 0 2
481 1023
476 1023
0 1 19 0 0 8320 0 0 41 41 0 3
198 797
198 1005
476 1005
2 0 20 0 0 4096 0 42 0 0 36 2
471 879
457 879
0 2 20 0 0 16384 0 0 42 40 0 5
264 938
264 954
335 954
335 879
471 879
1 1 17 0 0 4224 0 21 42 0 0 2
131 861
471 861
2 2 21 0 0 4224 0 44 43 0 0 3
311 933
311 760
475 760
2 1 22 0 0 12416 0 45 43 0 0 4
300 793
306 793
306 742
475 742
1 1 20 0 0 4224 0 20 44 0 0 3
133 938
275 938
275 933
1 1 19 0 0 0 0 22 45 0 0 3
133 797
264 797
264 793
1 4 23 0 0 4224 0 46 47 0 0 3
677 488
677 487
678 487
4 3 24 0 0 4224 0 51 47 0 0 4
461 593
624 593
624 496
632 496
4 2 25 0 0 4224 0 50 47 0 0 4
460 449
619 449
619 487
633 487
4 1 26 0 0 4224 0 49 47 0 0 4
454 354
624 354
624 478
632 478
0 3 27 0 0 4224 0 0 49 57 0 3
259 626
259 363
409 363
0 2 28 0 0 4096 0 0 49 52 0 3
377 449
377 354
409 354
2 1 29 0 0 4224 0 48 49 0 0 4
348 348
401 348
401 345
409 345
0 1 30 0 0 4096 0 0 48 53 0 3
243 417
243 348
312 348
0 0 31 0 0 4096 0 0 0 51 56 2
386 595
386 620
0 3 31 0 0 4224 0 0 50 0 0 3
386 616
386 458
415 458
0 2 28 0 0 0 0 0 50 54 0 3
359 471
359 449
415 449
1 1 30 0 0 4224 0 24 50 0 0 4
131 417
407 417
407 440
415 440
2 1 28 0 0 8320 0 54 51 0 0 4
341 471
403 471
403 584
416 584
2 2 32 0 0 4224 0 53 51 0 0 4
336 542
408 542
408 593
416 593
2 3 31 0 0 0 0 52 51 0 0 4
341 620
408 620
408 602
416 602
1 1 27 0 0 0 0 23 52 0 0 4
132 626
297 626
297 620
305 620
1 1 33 0 0 4224 0 26 53 0 0 4
131 558
292 558
292 542
300 542
1 1 34 0 0 4224 0 25 54 0 0 4
129 481
297 481
297 471
305 471
1 4 35 0 0 4224 0 55 57 0 0 2
313 185
313 184
1 3 36 0 0 4224 0 27 57 0 0 4
131 281
255 281
255 193
268 193
1 2 37 0 0 4224 0 28 57 0 0 4
129 204
260 204
260 184
268 184
2 1 38 0 0 4224 0 56 57 0 0 4
214 145
260 145
260 175
268 175
1 1 39 0 0 4224 0 29 56 0 0 4
131 140
170 140
170 145
178 145
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
70 49 175 74
88 57 156 72
9 Pagina 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
33 711 113 753
40 713 105 743
9 Pagina 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
29 1132 107 1174
35 1135 100 1165
9 Pagina 17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
56 1863 136 1905
63 1865 128 1895
9 Pagina 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 29
44 1888 268 1911
50 1891 261 1906
29 Aplicando a �lgebra booleana:
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 38
46 1967 226 2009
52 1969 219 1999
38 = (AB)' . ((A + B)')' =
(AB)' . (A+B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 39
51 1921 209 1963
57 1924 202 1954
39 F = ((AB) + A'B')' = 
(AB)' . (A'.B')'
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
