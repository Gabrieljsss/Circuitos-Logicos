CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
20 0 30 100 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 505 58 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4375 0 0
2
43401.3 0
0
13 Logic Switch~
5 245 56 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3616 0 0
2
43401.3 2
0
13 Logic Switch~
5 326 53 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7808 0 0
2
43401.3 1
0
13 Logic Switch~
5 406 59 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7498 0 0
2
43401.3 0
0
13 Logic Switch~
5 129 417 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9736 0 0
2
43401.3 0
0
14 Logic Display~
6 961 299 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9454 0 0
2
43401.3 0
0
14 Logic Display~
6 769 303 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4639 0 0
2
43401.3 0
0
14 Logic Display~
6 591 311 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3831 0 0
2
43401.3 0
0
14 Logic Display~
6 377 306 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3538 0 0
2
43401.3 0
0
4 4585
219 954 127 0 14 29
0 12 11 10 9 7 6 5 4 14
15 16 17 8 18
0
0 0 4848 0
4 4585
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
5949 0 0
2
43401.3 0
0
7 Ground~
168 206 255 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7130 0 0
2
43401.3 0
0
5 4013~
219 848 375 0 6 22
0 2 3 6 8 19 7
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U2A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 6 0
1 U
4115 0 0
2
43401.3 0
0
5 4013~
219 649 377 0 6 22
0 2 3 5 8 20 6
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
3197 0 0
2
43401.3 0
0
5 4013~
219 469 378 0 6 22
0 2 3 4 8 21 5
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U1A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
813 0 0
2
43401.3 0
0
5 4013~
219 273 387 0 6 22
0 2 3 13 8 22 4
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U6B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 4 0
1 U
3396 0 0
2
43401.3 2
0
7 Pulser~
4 166 613 0 10 12
0 23 24 25 26 0 0 5 5 3
7
0
0 0 4656 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6348 0 0
2
43401 0
0
28
5 2 0 0 0 0 0 12 12 0 0 4
878 357
878 303
824 303
824 339
5 2 0 0 0 0 0 13 13 0 0 5
679 359
689 359
689 308
625 308
625 341
5 2 0 0 0 0 0 14 14 0 0 5
499 360
512 360
512 306
445 306
445 342
5 2 0 0 0 0 0 15 15 0 0 5
303 369
315 369
315 317
249 317
249 351
0 1 4 0 0 8192 0 0 9 28 0 3
376 351
377 351
377 324
0 1 5 0 0 4096 0 0 8 27 0 2
591 359
591 329
0 1 6 0 0 4096 0 0 7 26 0 2
769 341
769 321
0 1 7 0 0 8192 0 0 6 16 0 3
909 316
909 317
961 317
0 4 8 0 0 8192 0 0 15 10 0 4
485 413
485 436
273 436
273 393
0 4 8 0 0 0 0 0 14 11 0 4
668 402
668 413
469 413
469 384
0 4 8 0 0 8192 0 0 13 12 0 4
887 381
887 402
649 402
649 383
13 4 8 0 0 8320 0 10 12 0 0 4
986 136
1019 136
1019 381
848 381
0 8 4 0 0 8320 0 0 10 28 0 3
338 351
338 154
922 154
0 7 5 0 0 8320 0 0 10 27 0 3
551 342
551 145
922 145
0 6 6 0 0 8320 0 0 10 26 0 3
714 341
714 136
922 136
6 5 7 0 0 8320 0 12 10 0 0 4
872 339
909 339
909 127
922 127
1 4 9 0 0 8320 0 2 10 0 0 3
257 56
257 118
922 118
1 3 10 0 0 8320 0 3 10 0 0 3
338 53
338 109
922 109
1 2 11 0 0 8320 0 4 10 0 0 3
418 59
418 100
922 100
1 1 12 0 0 4224 0 1 10 0 0 4
517 58
916 58
916 91
922 91
0 1 2 0 0 4224 0 0 12 22 0 3
649 249
848 249
848 318
0 1 2 0 0 0 0 0 13 23 0 3
469 249
649 249
649 320
0 1 2 0 0 0 0 0 14 24 0 3
272 249
469 249
469 321
1 1 2 0 0 0 0 11 15 0 0 3
206 249
273 249
273 330
1 3 13 0 0 12416 0 5 15 0 0 4
141 417
154 417
154 369
249 369
6 3 6 0 0 0 0 13 12 0 0 4
673 341
782 341
782 357
824 357
6 3 5 0 0 0 0 14 13 0 0 4
493 342
575 342
575 359
625 359
6 3 4 0 0 0 0 15 14 0 0 4
297 351
389 351
389 360
445 360
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
43 27 123 66
49 29 116 59
9 Pagina 15
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
