CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 2710 30 120 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 202 335 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7973 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 208 163 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8324 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 208 91 0 1 11
0 15
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
30 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 205 30 0 1 11
0 16
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3392 0 0
2
5.89862e-315 5.32571e-315
0
7 Ground~
168 611 378 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5283 0 0
2
5.89862e-315 0
0
7 Ground~
168 606 262 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6296 0 0
2
5.89862e-315 0
0
7 Ground~
168 759 153 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3981 0 0
2
5.89862e-315 0
0
7 Ground~
168 434 107 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7721 0 0
2
5.89862e-315 0
0
4 LED~
171 610 365 0 2 2
10 3 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D5
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3956 0 0
2
5.89862e-315 0
0
4 LED~
171 566 173 0 2 2
10 11 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3416 0 0
2
5.89862e-315 0
0
4 LED~
171 759 138 0 2 2
10 16 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8631 0 0
2
5.89862e-315 0
0
4 LED~
171 434 92 0 2 2
10 4 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3262 0 0
2
5.89862e-315 0
0
5 4049~
219 249 428 0 2 22
0 7 6
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 13 0
1 U
7874 0 0
2
5.89862e-315 5.34643e-315
0
8 2-In OR~
219 482 353 0 3 22
0 9 5 3
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 RpD
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
9834 0 0
2
5.89862e-315 5.3568e-315
0
5 4081~
219 328 417 0 3 22
0 8 6 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
4124 0 0
2
5.89862e-315 5.36716e-315
0
5 4081~
219 332 294 0 3 22
0 10 7 9
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
616 0 0
2
5.89862e-315 5.37752e-315
0
8 2-In OR~
219 478 167 0 3 22
0 13 12 11
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 RpC
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
799 0 0
2
43359.6 4
0
5 4081~
219 379 217 0 3 22
0 14 8 12
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
8849 0 0
2
43359.6 5
0
5 4049~
219 299 219 0 2 22
0 15 14
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 13 0
1 U
3871 0 0
2
43359.6 6
0
5 4049~
219 265 164 0 2 22
0 8 10
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 13 0
1 U
7991 0 0
2
43359.6 7
0
5 4081~
219 341 156 0 3 22
0 15 10 13
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
9107 0 0
2
43359.6 8
0
8 2-In OR~
219 348 82 0 3 22
0 16 15 4
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 RpB
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
7555 0 0
2
43359.6 9
0
26
1 2 2 0 0 4096 0 5 9 0 0 3
611 372
611 375
610 375
1 2 2 0 0 4224 0 6 10 0 0 4
606 256
606 212
566 212
566 183
1 2 2 0 0 0 0 7 11 0 0 2
759 147
759 148
1 2 2 0 0 0 0 8 12 0 0 2
434 101
434 102
1 0 3 0 0 4096 0 9 0 0 7 2
610 355
610 353
3 1 4 0 0 4224 0 22 12 0 0 2
381 82
434 82
3 0 3 0 0 4224 0 14 0 0 0 3
515 353
611 353
611 358
3 2 5 0 0 4224 0 15 14 0 0 3
349 417
469 417
469 362
2 2 6 0 0 8320 0 13 15 0 0 3
270 428
270 426
304 426
0 1 7 0 0 4096 0 0 13 13 0 3
219 335
219 428
234 428
0 1 8 0 0 4224 0 0 15 22 0 3
227 164
227 408
304 408
3 1 9 0 0 4224 0 16 14 0 0 3
353 294
469 294
469 344
1 2 7 0 0 4224 0 1 16 0 0 3
214 335
308 335
308 303
0 1 10 0 0 8320 0 0 16 21 0 3
307 165
308 165
308 285
3 1 11 0 0 12416 0 17 10 0 0 4
511 167
526 167
526 163
566 163
3 2 12 0 0 4224 0 18 17 0 0 3
400 217
465 217
465 176
3 1 13 0 0 8320 0 21 17 0 0 3
362 156
362 158
465 158
0 2 8 0 0 0 0 0 18 22 0 3
239 164
239 226
355 226
2 1 14 0 0 4224 0 19 18 0 0 3
320 219
355 219
355 208
0 1 15 0 0 8320 0 0 19 24 0 3
285 91
284 91
284 219
2 2 10 0 0 0 0 20 21 0 0 3
286 164
286 165
317 165
1 1 8 0 0 0 0 2 20 0 0 3
220 163
220 164
250 164
0 1 15 0 0 0 0 0 21 24 0 3
309 91
309 147
317 147
1 2 15 0 0 0 0 3 22 0 0 2
220 91
335 91
0 1 16 0 0 4096 0 0 22 26 0 3
328 30
328 73
335 73
1 1 16 0 0 4224 0 4 11 0 0 4
217 30
758 30
758 128
759 128
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
173 147 193 168
179 150 186 165
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
176 76 196 97
182 78 189 93
1 b
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
167 17 185 56
172 19 179 49
1 a
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
172 323 190 344
177 326 184 341
1 d
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
