CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 2190 30 120 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
31
13 Logic Switch~
5 801 464 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9828 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 718 470 0 1 11
0 19
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5906 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 620 473 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7780 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 443 488 0 1 11
0 5
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3518 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 309 475 0 1 11
0 18
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4262 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 176 485 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3944 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 267 76 0 1 11
0 30
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7617 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 180 79 0 1 11
0 27
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3202 0 0
2
5.89862e-315 0
0
7 Ground~
168 1301 635 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3969 0 0
2
5.89862e-315 0
0
4 LED~
171 1302 621 0 2 2
10 9 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9134 0 0
2
5.89862e-315 0
0
9 3-In AND~
219 1282 612 0 4 22
0 12 11 10 9
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 17 0
1 U
3615 0 0
2
5.89862e-315 0
0
5 4049~
219 1024 708 0 2 22
0 15 16
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 15 0
1 U
8504 0 0
2
5.89862e-315 5.34643e-315
0
5 4049~
219 1011 740 0 2 22
0 14 6
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 15 0
1 U
9765 0 0
2
5.89862e-315 5.32571e-315
0
5 4081~
219 1073 727 0 3 22
0 16 6 3
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 16 0
1 U
7195 0 0
2
5.89862e-315 5.30499e-315
0
5 4071~
219 1136 736 0 3 22
0 3 13 10
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 14 0
1 U
3832 0 0
2
5.89862e-315 5.26354e-315
0
5 4081~
219 1075 783 0 3 22
0 15 14 13
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 16 0
1 U
6663 0 0
2
5.89862e-315 0
0
5 4049~
219 1005 590 0 2 22
0 19 20
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 15 0
1 U
6215 0 0
2
5.89862e-315 5.34643e-315
0
5 4049~
219 1001 624 0 2 22
0 18 8
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 15 0
1 U
755 0 0
2
5.89862e-315 5.32571e-315
0
5 4081~
219 1054 609 0 3 22
0 20 8 4
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 16 0
1 U
9368 0 0
2
5.89862e-315 5.30499e-315
0
5 4071~
219 1117 618 0 3 22
0 4 17 11
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
3125 0 0
2
5.89862e-315 5.26354e-315
0
5 4081~
219 1056 665 0 3 22
0 18 19 17
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 16 0
1 U
3933 0 0
2
5.89862e-315 0
0
5 4081~
219 1066 545 0 3 22
0 22 5 21
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 13 0
1 U
3767 0 0
2
5.89862e-315 0
0
5 4071~
219 1127 498 0 3 22
0 23 21 12
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
3903 0 0
2
5.89862e-315 0
0
5 4081~
219 1064 489 0 3 22
0 24 7 23
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 13 0
1 U
9506 0 0
2
5.89862e-315 0
0
5 4049~
219 1004 502 0 2 22
0 5 7
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 15 0
1 U
4384 0 0
2
5.89862e-315 0
0
5 4049~
219 1015 470 0 2 22
0 22 24
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 15 0
1 U
9933 0 0
2
5.89862e-315 0
0
5 4071~
219 407 172 0 3 22
0 26 25 32
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 14 0
1 U
3754 0 0
2
5.89862e-315 0
0
5 4081~
219 310 123 0 3 22
0 30 27 26
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 13 0
1 U
973 0 0
2
5.89862e-315 0
0
5 4081~
219 312 244 0 3 22
0 29 28 25
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
3572 0 0
2
5.89862e-315 0
0
5 4069~
219 220 224 0 2 22
0 27 29
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U1B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
9628 0 0
2
5.89862e-315 0
0
5 4069~
219 222 276 0 2 22
0 30 33
0
0 0 608 0
4 4069
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 512 6 1 11 0
1 U
6617 0 0
2
5.89862e-315 0
0
43
0 1 3 0 0 4096 0 0 15 16 0 2
1117 727
1123 727
3 1 4 0 0 4224 0 19 20 0 0 2
1075 609
1104 609
3 0 4 0 0 0 0 19 0 0 22 2
1075 609
1096 609
2 0 5 0 0 4096 0 22 0 0 25 2
1042 554
1034 554
2 2 6 0 0 4224 0 13 14 0 0 3
1032 740
1049 740
1049 736
2 0 7 0 0 8320 0 25 0 0 28 3
1025 502
1025 503
1035 503
2 2 8 0 0 4224 0 18 19 0 0 3
1022 624
1030 624
1030 618
1 2 2 0 0 4224 0 9 10 0 0 3
1301 629
1301 631
1302 631
1 4 9 0 0 4224 0 10 11 0 0 3
1302 611
1302 612
1303 612
3 3 10 0 0 8320 0 15 11 0 0 3
1169 736
1258 736
1258 621
3 2 11 0 0 4224 0 20 11 0 0 4
1150 618
1234 618
1234 612
1258 612
3 1 12 0 0 8320 0 23 11 0 0 3
1160 498
1258 498
1258 603
3 2 13 0 0 8320 0 16 15 0 0 3
1096 783
1123 783
1123 745
0 2 14 0 0 8192 0 0 16 35 0 3
928 751
928 792
1051 792
0 1 15 0 0 8192 0 0 16 34 0 3
981 733
981 774
1051 774
3 1 3 0 0 4224 0 14 15 0 0 2
1094 727
1123 727
2 1 16 0 0 8320 0 12 14 0 0 3
1045 708
1049 708
1049 718
0 1 14 0 0 0 0 0 13 35 0 3
961 751
996 751
996 740
3 2 17 0 0 4224 0 21 20 0 0 3
1077 665
1077 627
1104 627
0 1 18 0 0 8192 0 0 21 33 0 3
970 645
970 656
1032 656
0 2 19 0 0 8192 0 0 21 32 0 3
943 627
943 674
1032 674
0 1 4 0 0 0 0 0 20 0 0 3
1078 610
1078 609
1104 609
2 1 20 0 0 8320 0 17 19 0 0 3
1026 590
1030 590
1030 600
3 2 21 0 0 8320 0 22 23 0 0 3
1087 545
1114 545
1114 507
0 2 5 0 0 4096 0 0 22 31 0 4
981 546
1034 546
1034 554
1042 554
0 1 22 0 0 4096 0 0 22 30 0 3
957 524
1042 524
1042 536
3 1 23 0 0 4224 0 24 23 0 0 2
1085 489
1114 489
0 2 7 0 0 0 0 0 24 0 0 3
1031 503
1040 503
1040 498
2 1 24 0 0 8320 0 26 24 0 0 3
1036 470
1040 470
1040 480
1 1 22 0 0 8320 0 1 26 0 0 5
813 464
813 532
957 532
957 470
1000 470
1 1 5 0 0 8320 0 4 25 0 0 5
455 488
455 550
981 550
981 502
989 502
1 1 19 0 0 8320 0 2 17 0 0 5
730 470
730 627
967 627
967 590
990 590
1 1 18 0 0 8320 0 5 18 0 0 4
321 475
321 645
986 645
986 624
1 1 15 0 0 8320 0 3 12 0 0 5
632 473
632 733
996 733
996 708
1009 708
1 0 14 0 0 8320 0 6 0 0 0 3
188 485
188 751
970 751
3 2 25 0 0 8320 0 29 27 0 0 3
333 244
394 244
394 181
3 1 26 0 0 4224 0 28 27 0 0 3
331 123
394 123
394 163
0 2 27 0 0 4096 0 0 28 43 0 2
192 132
286 132
0 2 28 0 0 4224 0 0 29 0 0 3
236 275
288 275
288 253
2 1 29 0 0 4224 0 30 29 0 0 3
241 224
288 224
288 235
0 1 30 0 0 8320 0 0 31 42 0 4
279 93
166 93
166 276
207 276
1 1 30 0 0 0 0 7 28 0 0 3
279 76
279 114
286 114
1 1 27 0 0 4224 0 8 30 0 0 3
192 79
192 224
205 224
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
61 22 79 43
66 25 73 40
1 c
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
233 407 358 446
239 409 351 439
15 Primeiro numero
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
674 402 792 441
680 405 785 435
14 Segundo numero
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
118 448 153 469
124 451 146 466
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
568 447 603 468
574 450 596 465
3 MSB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
