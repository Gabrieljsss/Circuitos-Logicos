CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 50 30 140 10
176 86 1918 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 182 457 279
42991634 0
0
6 Title:
5 Name:
0
0
0
26
13 Logic Switch~
5 896 289 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -13 12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6118 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 139 579 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
5.89871e-315 5.26354e-315
0
13 Logic Switch~
5 138 620 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6357 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 139 548 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
319 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 140 507 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3976 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 483 424 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7634 0 0
2
43434.5 0
0
13 Logic Switch~
5 196 297 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
523 0 0
2
43434.5 1
0
13 Logic Switch~
5 202 133 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6748 0 0
2
43434.5 2
0
13 Logic Switch~
5 149 187 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -13 8 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6901 0 0
2
5.89871e-315 0
0
5 4071~
219 1001 375 0 3 22
0 6 7 2
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U7A
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
842 0 0
2
5.89871e-315 0
0
5 4071~
219 933 376 0 3 22
0 8 9 3
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U3D
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
3277 0 0
2
5.89871e-315 0
0
5 4071~
219 870 377 0 3 22
0 11 10 4
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U3C
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
4212 0 0
2
5.89871e-315 0
0
5 4081~
219 236 609 0 3 22
0 12 13 6
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
4720 0 0
2
5.89871e-315 0
0
5 4081~
219 233 569 0 3 22
0 12 14 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
5551 0 0
2
5.89871e-315 0
0
5 4081~
219 234 532 0 3 22
0 12 15 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
6986 0 0
2
5.89871e-315 0
0
5 4049~
219 755 129 0 2 22
0 10 18
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5B
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
8745 0 0
2
43434.5 3
0
5 4081~
219 722 138 0 3 22
0 18 17 16
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
9592 0 0
2
43434.5 4
0
5 4071~
219 566 126 0 3 22
0 10 21 20
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
8748 0 0
2
43434.5 5
0
5 4049~
219 324 300 0 2 22
0 17 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
7168 0 0
2
43434.5 6
0
5 4081~
219 492 107 0 3 22
0 9 21 23
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
631 0 0
2
43434.5 7
0
5 4071~
219 348 96 0 3 22
0 7 23 22
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9466 0 0
2
43434.5 8
0
12 Hex Display~
7 956 230 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3266 0 0
2
43434.5 9
0
7 Pulser~
4 150 91 0 10 12
0 26 27 28 29 0 0 5 5 2
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7693 0 0
2
5.89871e-315 5.26354e-315
0
5 4027~
219 804 241 0 7 32
0 25 16 24 19 12 30 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3723 0 0
2
5.89871e-315 5.30499e-315
0
5 4027~
219 603 239 0 7 32
0 25 19 24 20 12 31 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3440 0 0
2
5.89871e-315 5.32571e-315
0
5 4027~
219 408 238 0 7 32
0 25 22 24 9 12 32 10
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6263 0 0
2
5.89871e-315 5.34643e-315
0
41
3 1 2 0 0 4224 0 10 22 0 0 4
1004 345
1004 272
965 272
965 254
3 2 3 0 0 12416 0 11 22 0 0 4
936 346
936 319
959 319
959 254
3 3 4 0 0 8320 0 12 22 0 0 4
873 347
873 310
953 310
953 254
1 4 5 0 0 8320 0 1 22 0 0 3
908 289
908 254
947 254
3 1 6 0 0 4224 0 13 10 0 0 3
257 609
995 609
995 391
0 2 7 0 0 4096 0 0 10 31 0 4
828 139
1085 139
1085 391
1013 391
3 1 8 0 0 4224 0 14 11 0 0 3
254 569
927 569
927 392
0 2 9 0 0 8320 0 0 11 29 0 4
635 277
635 429
945 429
945 392
0 2 10 0 0 12416 0 0 12 21 0 5
432 152
456 152
456 470
882 470
882 393
3 1 11 0 0 4224 0 15 12 0 0 3
255 532
864 532
864 393
0 1 12 0 0 4096 0 0 13 14 0 3
194 560
194 600
212 600
1 2 13 0 0 8320 0 3 13 0 0 3
150 620
150 618
212 618
1 2 14 0 0 8320 0 2 14 0 0 3
151 579
151 578
209 578
0 1 12 0 0 4096 0 0 14 19 0 3
176 507
176 560
209 560
1 2 15 0 0 8320 0 4 15 0 0 3
151 548
151 541
210 541
0 1 12 0 0 0 0 0 15 19 0 3
203 507
203 523
210 523
0 5 12 0 0 8192 0 0 24 18 0 3
602 507
804 507
804 247
0 5 12 0 0 8192 0 0 25 19 0 3
408 507
603 507
603 245
1 5 12 0 0 8320 0 5 26 0 0 3
152 507
408 507
408 244
0 1 10 0 0 0 0 0 16 21 0 4
531 121
531 41
776 41
776 129
7 1 10 0 0 0 0 26 18 0 0 4
432 202
432 121
585 121
585 117
3 2 16 0 0 8320 0 17 24 0 0 3
697 138
697 205
780 205
0 2 17 0 0 8320 0 0 17 35 0 4
278 300
278 319
742 319
742 147
2 1 18 0 0 4224 0 16 17 0 0 2
740 129
742 129
0 4 19 0 0 4224 0 0 24 28 0 3
529 355
780 355
780 223
3 4 20 0 0 4224 0 18 25 0 0 3
539 126
539 221
579 221
0 2 21 0 0 4096 0 0 18 34 0 3
512 147
585 147
585 135
1 2 19 0 0 0 0 6 25 0 0 4
495 424
529 424
529 203
579 203
0 4 9 0 0 0 0 0 26 33 0 5
627 195
642 195
642 277
384 277
384 220
3 2 22 0 0 4224 0 21 26 0 0 3
321 96
321 202
384 202
7 1 7 0 0 8320 0 24 21 0 0 3
828 205
828 87
367 87
3 2 23 0 0 8320 0 20 21 0 0 3
467 107
467 105
367 105
7 1 9 0 0 0 0 25 20 0 0 3
627 203
627 98
512 98
2 2 21 0 0 8320 0 19 20 0 0 3
345 300
512 300
512 116
1 1 17 0 0 0 0 7 19 0 0 3
208 297
208 300
309 300
3 3 24 0 0 8320 0 25 24 0 0 3
579 212
579 214
780 214
3 3 24 0 0 0 0 26 25 0 0 3
384 211
384 212
579 212
1 3 24 0 0 0 0 8 26 0 0 3
214 133
214 211
384 211
1 1 25 0 0 8192 0 25 24 0 0 3
603 182
603 184
804 184
1 1 25 0 0 0 0 26 25 0 0 3
408 181
408 182
603 182
1 1 25 0 0 4224 0 9 26 0 0 4
161 187
367 187
367 181
408 181
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
122 340 274 364
127 342 268 358
18 1 = multiplos de 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
121 319 273 343
126 321 267 337
18 0 = multiplos de 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
130 285 173 309
132 287 170 303
5 Input
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
142 121 189 145
146 123 184 139
5 Clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
802 153 819 177
806 154 814 170
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
591 142 610 166
596 144 604 160
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
397 140 414 164
401 142 409 158
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
89 177 127 199
96 180 119 196
3 gnd
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
49 492 103 516
53 494 98 510
6 Ativar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
46 523 80 547
51 524 74 540
3 MSB
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
