CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
1070 260 30 80 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
71
13 Logic Switch~
5 925 213 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3280 0 0
2
5.89867e-315 0
0
13 Logic Switch~
5 817 213 0 1 11
0 63
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3122 0 0
2
5.89867e-315 5.26354e-315
0
13 Logic Switch~
5 724 202 0 1 11
0 62
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6242 0 0
2
5.89867e-315 5.30499e-315
0
13 Logic Switch~
5 620 202 0 1 11
0 60
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8862 0 0
2
5.89867e-315 5.32571e-315
0
13 Logic Switch~
5 552 199 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3202 0 0
2
5.89867e-315 5.34643e-315
0
13 Logic Switch~
5 46 195 0 10 11
0 51 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5657 0 0
2
5.89867e-315 5.3568e-315
0
13 Logic Switch~
5 135 194 0 1 11
0 52
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3554 0 0
2
5.89867e-315 5.36716e-315
0
13 Logic Switch~
5 239 194 0 1 11
0 53
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4316 0 0
2
5.89867e-315 5.37752e-315
0
13 Logic Switch~
5 332 205 0 10 11
0 54 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3739 0 0
2
5.89867e-315 5.38788e-315
0
13 Logic Switch~
5 440 205 0 1 11
0 55
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7606 0 0
2
5.89867e-315 5.39306e-315
0
14 Logic Display~
6 3040 1390 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
43403.4 0
0
14 Logic Display~
6 3032 1280 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
369 0 0
2
43403.4 1
0
14 Logic Display~
6 3029 1080 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8773 0 0
2
43403.4 2
0
14 Logic Display~
6 3031 771 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7981 0 0
2
43403.4 3
0
8 2-In OR~
219 2526 1329 0 3 22
0 10 9 3
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 33 0
1 U
4205 0 0
2
43403.4 4
0
9 2-In AND~
219 2491 1370 0 3 22
0 11 6 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 34 0
1 U
3375 0 0
2
43403.4 5
0
5 4030~
219 2432 1357 0 3 22
0 12 12 11
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 35 0
1 U
719 0 0
2
43403.4 6
0
9 2-In AND~
219 2415 1296 0 3 22
0 13 12 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 34 0
1 U
3749 0 0
2
43403.4 7
0
5 4049~
219 2364 1285 0 2 22
0 6 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 29 0
1 U
3871 0 0
2
43403.4 8
0
8 2-In OR~
219 2770 1131 0 3 22
0 15 14 4
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 33 0
1 U
4393 0 0
2
43403.4 9
0
9 2-In AND~
219 2714 1222 0 3 22
0 16 6 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
6229 0 0
2
43403.4 10
0
8 2-In OR~
219 2641 1182 0 3 22
0 18 17 16
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
3757 0 0
2
43403.4 11
0
8 2-In OR~
219 2544 1144 0 3 22
0 20 19 18
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
352 0 0
2
43403.4 12
0
9 2-In AND~
219 2483 1112 0 3 22
0 7 21 20
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
3372 0 0
2
43403.4 13
0
9 2-In AND~
219 2411 1115 0 3 22
0 23 22 21
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
4911 0 0
2
43403.4 14
0
9 2-In AND~
219 2478 1172 0 3 22
0 24 12 19
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
7574 0 0
2
43403.4 15
0
9 2-In AND~
219 2478 1222 0 3 22
0 24 8 17
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
6601 0 0
2
43403.4 16
0
5 4049~
219 2359 1164 0 2 22
0 7 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 29 0
1 U
8531 0 0
2
43403.4 17
0
5 4049~
219 2359 1124 0 2 22
0 8 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 29 0
1 U
6532 0 0
2
43403.4 18
0
5 4049~
219 2359 1105 0 2 22
0 12 23
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 29 0
1 U
3621 0 0
2
43403.4 19
0
9 2-In AND~
219 2410 1029 0 3 22
0 25 7 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
5174 0 0
2
43403.4 20
0
5 4049~
219 2353 1017 0 2 22
0 6 25
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 29 0
1 U
5452 0 0
2
43403.4 21
0
8 2-In OR~
219 2953 804 0 3 22
0 27 26 5
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 31 0
1 U
3626 0 0
2
43403.4 22
0
9 2-In AND~
219 2896 909 0 3 22
0 28 6 26
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
3806 0 0
2
43403.4 23
0
8 2-In OR~
219 2791 849 0 3 22
0 30 29 28
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
3389 0 0
2
43403.4 24
0
8 2-In OR~
219 2679 881 0 3 22
0 32 31 29
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
9156 0 0
2
43403.4 25
0
8 2-In OR~
219 2679 774 0 3 22
0 34 33 30
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
5810 0 0
2
43403.4 26
0
9 2-In AND~
219 2622 924 0 3 22
0 36 35 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
8260 0 0
2
43403.4 27
0
9 2-In AND~
219 2570 958 0 3 22
0 37 40 35
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
7286 0 0
2
43403.4 28
0
9 2-In AND~
219 2568 905 0 3 22
0 38 39 36
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
3689 0 0
2
43403.4 29
0
5 4049~
219 2509 945 0 2 22
0 8 37
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 29 0
1 U
4485 0 0
2
43403.4 30
0
5 4049~
219 2511 917 0 2 22
0 12 39
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 23 0
1 U
4370 0 0
2
43403.4 31
0
5 4049~
219 2509 894 0 2 22
0 7 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 23 0
1 U
7483 0 0
2
43403.4 32
0
9 2-In AND~
219 2513 846 0 3 22
0 41 8 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
4214 0 0
2
43403.4 33
0
9 2-In AND~
219 2514 798 0 3 22
0 41 12 33
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
9254 0 0
2
43403.4 34
0
9 2-In AND~
219 2515 741 0 3 22
0 41 7 34
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
7515 0 0
2
43403.4 35
0
5 4049~
219 2382 727 0 2 22
0 40 41
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 23 0
1 U
9241 0 0
2
43403.4 36
0
9 2-In AND~
219 2434 672 0 3 22
0 42 40 27
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
3783 0 0
2
43403.4 37
0
5 4049~
219 2382 654 0 2 22
0 6 42
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 23 0
1 U
5226 0 0
2
43403.4 38
0
9 2-In AND~
219 2592 518 0 3 22
0 6 44 43
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
6496 0 0
2
43403.4 39
0
8 2-In OR~
219 2512 568 0 3 22
0 46 45 44
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
6819 0 0
2
43403.4 40
0
8 2-In OR~
219 2430 588 0 3 22
0 12 8 45
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U18D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
6832 0 0
2
43403.4 41
0
8 2-In OR~
219 2431 551 0 3 22
0 40 7 46
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U18C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
7222 0 0
2
43403.4 42
0
14 Logic Display~
6 1742 922 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4676 0 0
2
5.89867e-315 5.39824e-315
0
14 Logic Display~
6 1736 855 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9334 0 0
2
5.89867e-315 5.40342e-315
0
14 Logic Display~
6 1729 777 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4758 0 0
2
5.89867e-315 5.4086e-315
0
14 Logic Display~
6 1728 711 0 1 2
10 40
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6695 0 0
2
5.89867e-315 5.41378e-315
0
14 Logic Display~
6 1907 1159 0 1 2
10 48
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8212 0 0
2
5.89867e-315 5.41896e-315
0
5 4069~
219 1565 1206 0 2 22
0 49 6
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
3922 0 0
2
5.89867e-315 5.42414e-315
0
6 74LS83
105 1775 1161 0 14 29
0 2 2 2 51 2 2 2 50 6
65 66 67 48 68
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
7610 0 0
2
5.89867e-315 5.42933e-315
0
7 Ground~
168 1224 903 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6131 0 0
2
5.89867e-315 5.43192e-315
0
6 74LS83
105 1505 832 0 14 29
0 58 57 56 47 52 53 54 55 2
40 7 12 8 49
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
7187 0 0
2
5.89867e-315 5.43451e-315
0
5 4030~
219 1143 452 0 3 22
0 47 63 56
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9198 0 0
2
5.89867e-315 5.4371e-315
0
5 4030~
219 1276 551 0 3 22
0 59 62 57
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
9468 0 0
2
5.89867e-315 5.43969e-315
0
5 4030~
219 1403 657 0 3 22
0 61 60 58
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
5160 0 0
2
5.89867e-315 5.44228e-315
0
5 4071~
219 1073 535 0 3 22
0 63 47 59
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
7647 0 0
2
5.89867e-315 5.44487e-315
0
5 4071~
219 1164 626 0 3 22
0 62 59 61
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7210 0 0
2
5.89867e-315 5.44746e-315
0
14 Logic Display~
6 1097 313 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7128 0 0
2
5.89867e-315 5.45005e-315
0
14 Logic Display~
6 1213 426 0 1 2
10 56
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5367 0 0
2
5.89867e-315 5.45264e-315
0
14 Logic Display~
6 1357 526 0 1 2
10 57
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7140 0 0
2
5.89867e-315 5.45523e-315
0
14 Logic Display~
6 1472 642 0 1 2
10 58
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4903 0 0
2
5.89867e-315 5.45782e-315
0
128
1 3 3 0 0 4224 0 12 15 0 0 4
3032 1298
2558 1298
2558 1329
2559 1329
1 3 4 0 0 8320 0 13 20 0 0 3
3029 1098
3029 1131
2803 1131
1 3 5 0 0 8320 0 14 33 0 0 3
3031 789
3031 804
2986 804
0 0 6 0 0 12288 0 0 0 89 77 5
1684 1206
1684 1044
2100 1044
2100 496
2131 496
1 0 7 0 0 8192 0 56 0 0 78 5
1729 795
1900 795
1900 388
2222 388
2222 490
0 0 8 0 0 8192 0 0 0 87 79 5
1740 946
2061 946
2061 453
2307 453
2307 486
0 1 8 0 0 12288 0 0 11 79 0 4
2307 1419
2330 1419
2330 1408
3040 1408
2 3 9 0 0 8320 0 15 16 0 0 3
2513 1338
2512 1338
2512 1370
1 3 10 0 0 8320 0 15 18 0 0 3
2513 1320
2513 1296
2436 1296
1 3 11 0 0 4224 0 16 17 0 0 3
2467 1361
2467 1357
2465 1357
0 2 6 0 0 0 0 0 16 77 0 3
2131 1385
2467 1385
2467 1379
2 0 12 0 0 4096 0 17 0 0 80 2
2416 1366
2271 1366
1 0 12 0 0 0 0 17 0 0 80 2
2416 1348
2271 1348
1 2 13 0 0 8320 0 18 19 0 0 3
2391 1287
2391 1285
2385 1285
0 2 12 0 0 0 0 0 18 80 0 3
2271 1308
2391 1308
2391 1305
0 1 6 0 0 0 0 0 19 77 0 3
2131 1286
2349 1286
2349 1285
2 3 14 0 0 4224 0 20 21 0 0 3
2757 1140
2757 1222
2735 1222
1 3 15 0 0 8320 0 20 31 0 0 3
2757 1122
2757 1029
2431 1029
1 3 16 0 0 4224 0 21 22 0 0 4
2690 1213
2690 1197
2674 1197
2674 1182
0 2 6 0 0 4096 0 0 21 77 0 3
2131 1255
2690 1255
2690 1231
2 3 17 0 0 4224 0 22 27 0 0 3
2628 1191
2499 1191
2499 1222
1 3 18 0 0 8320 0 22 23 0 0 3
2628 1173
2628 1144
2577 1144
2 3 19 0 0 8320 0 23 26 0 0 3
2531 1153
2531 1172
2499 1172
1 3 20 0 0 4224 0 23 24 0 0 3
2531 1135
2504 1135
2504 1112
3 2 21 0 0 8320 0 25 24 0 0 3
2432 1115
2432 1121
2459 1121
2 2 22 0 0 4224 0 25 29 0 0 2
2387 1124
2380 1124
1 2 23 0 0 8320 0 25 30 0 0 3
2387 1106
2387 1105
2380 1105
0 2 8 0 0 0 0 0 27 79 0 3
2307 1234
2454 1234
2454 1231
0 1 24 0 0 8192 0 0 27 30 0 3
2396 1164
2396 1213
2454 1213
2 1 24 0 0 4224 0 28 26 0 0 3
2380 1164
2454 1164
2454 1163
0 2 12 0 0 4096 0 0 26 80 0 3
2271 1184
2454 1184
2454 1181
0 1 7 0 0 0 0 0 28 78 0 2
2222 1164
2344 1164
0 1 8 0 0 0 0 0 29 79 0 2
2307 1124
2344 1124
0 1 12 0 0 0 0 0 30 80 0 2
2271 1105
2344 1105
0 1 7 0 0 0 0 0 24 78 0 3
2222 1089
2459 1089
2459 1103
1 2 25 0 0 4224 0 31 32 0 0 3
2386 1020
2374 1020
2374 1017
0 2 7 0 0 0 0 0 31 78 0 4
2222 1042
2237 1042
2237 1038
2386 1038
0 1 6 0 0 0 0 0 32 77 0 2
2131 1017
2338 1017
2 3 26 0 0 8320 0 33 34 0 0 3
2940 813
2917 813
2917 909
1 3 27 0 0 8320 0 33 48 0 0 3
2940 795
2940 672
2455 672
1 3 28 0 0 4224 0 34 35 0 0 3
2872 900
2872 849
2824 849
0 2 6 0 0 4096 0 0 34 77 0 3
2131 997
2872 997
2872 918
2 3 29 0 0 8320 0 35 36 0 0 3
2778 858
2778 881
2712 881
1 3 30 0 0 4224 0 35 37 0 0 3
2778 840
2712 840
2712 774
2 3 31 0 0 8320 0 36 38 0 0 3
2666 890
2643 890
2643 924
1 3 32 0 0 4224 0 36 44 0 0 4
2666 872
2549 872
2549 846
2534 846
2 3 33 0 0 4224 0 37 45 0 0 3
2666 783
2535 783
2535 798
1 3 34 0 0 8320 0 37 46 0 0 4
2666 765
2666 756
2536 756
2536 741
2 3 35 0 0 4224 0 38 39 0 0 3
2598 933
2598 958
2591 958
3 1 36 0 0 4224 0 40 38 0 0 3
2589 905
2589 915
2598 915
1 2 37 0 0 8320 0 39 41 0 0 3
2546 949
2546 945
2530 945
1 2 38 0 0 8320 0 40 43 0 0 3
2544 896
2544 894
2530 894
2 2 39 0 0 4224 0 40 42 0 0 3
2544 914
2532 914
2532 917
0 2 40 0 0 4096 0 0 39 81 0 3
2178 971
2546 971
2546 967
0 1 8 0 0 0 0 0 41 79 0 2
2307 945
2494 945
0 1 12 0 0 4096 0 0 42 80 0 2
2271 917
2496 917
0 1 7 0 0 0 0 0 43 78 0 2
2222 894
2494 894
0 2 8 0 0 0 0 0 44 79 0 2
2307 855
2489 855
0 1 41 0 0 4224 0 0 44 62 0 3
2443 727
2443 837
2489 837
0 2 12 0 0 0 0 0 45 80 0 3
2271 809
2490 809
2490 807
0 1 41 0 0 0 0 0 45 62 0 4
2416 727
2416 788
2490 788
2490 789
2 1 41 0 0 0 0 47 46 0 0 3
2403 727
2491 727
2491 732
0 2 7 0 0 0 0 0 46 78 0 3
2222 755
2491 755
2491 750
0 1 40 0 0 0 0 0 47 81 0 2
2178 727
2367 727
2 0 40 0 0 0 0 48 0 0 81 2
2410 681
2178 681
1 2 42 0 0 4224 0 48 49 0 0 3
2410 663
2410 654
2403 654
0 1 6 0 0 0 0 0 49 77 0 2
2131 654
2367 654
3 0 43 0 0 4224 0 50 0 0 0 2
2613 518
2648 518
1 0 6 0 0 0 0 50 0 0 77 2
2568 509
2131 509
2 3 44 0 0 8320 0 50 51 0 0 3
2568 527
2545 527
2545 568
2 3 45 0 0 8320 0 51 52 0 0 3
2499 577
2499 588
2463 588
1 3 46 0 0 8320 0 51 53 0 0 3
2499 559
2499 551
2464 551
2 0 8 0 0 0 0 52 0 0 79 2
2417 597
2307 597
1 0 12 0 0 0 0 52 0 0 80 2
2417 579
2271 579
2 0 7 0 0 0 0 53 0 0 78 2
2418 560
2222 560
1 0 40 0 0 0 0 53 0 0 81 2
2418 542
2178 542
0 0 6 0 0 8320 0 0 0 0 11 4
2136 490
2131 490
2131 1385
2155 1385
0 0 7 0 0 8320 0 0 0 0 0 3
2220 1176
2222 1176
2222 487
0 0 8 0 0 8320 0 0 0 0 7 4
2308 483
2307 483
2307 1419
2330 1419
1 0 12 0 0 16512 0 55 0 0 12 6
1736 873
1955 873
1955 423
2271 423
2271 1366
2294 1366
1 0 40 0 0 16512 0 57 0 0 54 6
1728 729
1863 729
1863 356
2178 356
2178 971
2196 971
0 0 47 0 0 8192 0 0 0 125 114 3
974 354
974 353
1035 353
0 1 2 0 0 4096 0 0 61 101 0 3
1280 885
1224 885
1224 897
10 1 40 0 0 0 0 62 57 0 0 6
1537 823
1594 823
1594 720
1697 720
1697 729
1728 729
0 1 7 0 0 0 0 0 56 0 0 3
1702 792
1702 795
1729 795
12 1 12 0 0 0 0 62 55 0 0 6
1537 841
1632 841
1632 862
1703 862
1703 873
1736 873
13 1 8 0 0 0 0 62 54 0 0 7
1537 850
1580 850
1580 937
1708 937
1708 946
1742 946
1742 940
13 1 48 0 0 8320 0 60 58 0 0 3
1807 1179
1807 1177
1907 1177
2 9 6 0 0 0 0 59 60 0 0 2
1586 1206
1743 1206
14 1 49 0 0 8320 0 62 59 0 0 4
1537 877
1544 877
1544 1206
1550 1206
0 8 50 0 0 8320 0 0 60 92 0 3
560 334
560 1188
1743 1188
1 0 50 0 0 0 0 5 0 0 0 3
564 199
560 199
560 349
1 4 51 0 0 8320 0 6 60 0 0 3
58 195
58 1152
1743 1152
0 7 2 0 0 8320 0 0 60 95 0 3
1454 1170
1454 1179
1743 1179
0 6 2 0 0 0 0 0 60 96 0 3
1454 1161
1454 1170
1743 1170
0 5 2 0 0 0 0 0 60 97 0 3
1454 1143
1454 1161
1743 1161
0 3 2 0 0 0 0 0 60 98 0 3
1454 1133
1454 1143
1743 1143
0 2 2 0 0 0 0 0 60 99 0 3
1454 1125
1454 1134
1743 1134
0 1 2 0 0 0 0 0 60 101 0 3
1454 885
1454 1125
1743 1125
11 0 7 0 0 0 0 62 0 0 85 5
1537 832
1608 832
1608 783
1705 783
1705 795
0 9 2 0 0 0 0 0 62 0 0 3
1264 885
1473 885
1473 877
1 5 52 0 0 8320 0 7 62 0 0 3
147 194
147 832
1473 832
1 6 53 0 0 8320 0 8 62 0 0 3
251 194
251 841
1473 841
1 7 54 0 0 8320 0 9 62 0 0 3
344 205
344 850
1473 850
1 8 55 0 0 8320 0 10 62 0 0 3
452 205
452 859
1473 859
0 4 47 0 0 4224 0 0 62 114 0 3
1060 353
1060 823
1473 823
0 3 56 0 0 4224 0 0 62 113 0 3
1186 452
1186 814
1473 814
0 2 57 0 0 4224 0 0 62 112 0 3
1331 551
1331 805
1473 805
0 1 58 0 0 4224 0 0 62 111 0 3
1441 660
1441 796
1473 796
0 3 59 0 0 4096 0 0 66 120 0 2
1113 535
1106 535
3 1 58 0 0 0 0 65 71 0 0 3
1436 657
1436 660
1472 660
3 1 57 0 0 0 0 64 70 0 0 3
1309 551
1357 551
1357 544
3 1 56 0 0 0 0 63 69 0 0 3
1176 452
1213 452
1213 444
0 1 47 0 0 0 0 0 68 0 0 3
1032 353
1097 353
1097 331
1 2 60 0 0 8320 0 4 65 0 0 3
632 202
632 666
1387 666
3 1 61 0 0 4224 0 67 65 0 0 4
1197 626
1323 626
1323 648
1387 648
0 2 59 0 0 4096 0 0 67 120 0 3
1117 535
1117 635
1151 635
0 1 62 0 0 8192 0 0 67 119 0 3
1023 560
1023 617
1151 617
1 2 62 0 0 8320 0 3 64 0 0 3
736 202
736 560
1260 560
0 1 59 0 0 4224 0 0 64 0 0 4
1109 535
1254 535
1254 542
1260 542
0 2 47 0 0 0 0 0 66 124 0 3
1048 443
1048 544
1060 544
0 1 63 0 0 8192 0 0 66 123 0 3
829 460
829 526
1060 526
1 2 63 0 0 8320 0 2 63 0 0 3
829 213
829 461
1127 461
0 1 47 0 0 0 0 0 63 0 0 3
1043 440
1043 443
1127 443
1 0 47 0 0 0 0 1 0 0 121 5
937 213
974 213
974 431
1048 431
1048 443
0 1 60 0 0 0 0 0 4 0 0 3
635 214
635 202
632 202
0 1 52 0 0 0 0 0 7 0 0 3
150 206
150 194
147 194
0 0 64 0 0 4224 0 0 0 0 0 2
128 1205
128 1188
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
3083 1371 3123 1394
3091 1375 3114 1390
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 27
3144 988 3366 1011
3153 991 3356 1006
27 SAIDAS QUE FORMAM A UNIDADE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1868 1086 2013 1109
1876 1090 2004 1105
17 Saida das dezenas
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2648 504 2670 528
2655 509 2662 525
1 E
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2810 1121 2832 1145
2817 1126 2824 1142
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2560 1313 2582 1337
2567 1319 2574 1335
1 H
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
2566 1412 2588 1436
2573 1417 2580 1433
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
72 108 150 129
77 111 144 126
9 questao 2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
