CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 390 16 60 10
176 86 1918 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 182 457 279
42991634 0
0
6 Title:
5 Name:
0
0
0
82
13 Logic Switch~
5 641 1798 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6421 0 0
2
5.8987e-315 0
0
13 Logic Switch~
5 647 1642 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7743 0 0
2
5.8987e-315 5.26354e-315
0
13 Logic Switch~
5 650 1585 0 10 11
0 29 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9840 0 0
2
5.8987e-315 5.30499e-315
0
13 Logic Switch~
5 649 1538 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6910 0 0
2
5.8987e-315 5.32571e-315
0
13 Logic Switch~
5 643 1728 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
449 0 0
2
5.8987e-315 5.34643e-315
0
13 Logic Switch~
5 641 1766 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8761 0 0
2
5.8987e-315 5.3568e-315
0
13 Logic Switch~
5 820 1707 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
5.8987e-315 5.36716e-315
0
13 Logic Switch~
5 647 1689 0 10 11
0 27 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7393 0 0
2
5.8987e-315 5.37752e-315
0
13 Logic Switch~
5 657 1246 0 1 11
0 44
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7699 0 0
2
5.8987e-315 5.38788e-315
0
13 Logic Switch~
5 321 471 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6638 0 0
2
43429.4 0
0
13 Logic Switch~
5 154 971 0 1 11
0 49
0
0 0 21360 0
2 0V
-10 -15 4 -7
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4595 0 0
2
43429.4 1
0
13 Logic Switch~
5 830 1264 0 1 11
0 59
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9395 0 0
2
5.8987e-315 5.39824e-315
0
13 Logic Switch~
5 651 1323 0 1 11
0 61
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3303 0 0
2
5.8987e-315 5.40342e-315
0
13 Logic Switch~
5 653 1285 0 10 11
0 62 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4498 0 0
2
5.8987e-315 5.4086e-315
0
13 Logic Switch~
5 659 1095 0 1 11
0 63
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9728 0 0
2
5.8987e-315 5.41378e-315
0
13 Logic Switch~
5 660 1142 0 1 11
0 64
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3789 0 0
2
5.8987e-315 5.41896e-315
0
13 Logic Switch~
5 657 1199 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3978 0 0
2
5.8987e-315 5.42414e-315
0
13 Logic Switch~
5 737 584 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3494 0 0
2
5.8987e-315 5.42933e-315
0
13 Logic Switch~
5 727 651 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3507 0 0
2
5.8987e-315 5.43192e-315
0
7 Pulser~
4 312 418 0 10 12
0 70 71 51 72 0 0 30 30 19
8
0
0 0 4656 0
0
3 V27
-11 -28 10 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5151 0 0
2
5.8987e-315 0
0
5 4049~
219 437 1204 0 2 22
0 2 3
0
0 0 624 512
4 4049
-7 -24 21 -16
4 U26B
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 24 0
1 U
3701 0 0
2
5.8987e-315 0
0
5 4049~
219 437 1096 0 2 22
0 7 8
0
0 0 624 512
4 4049
-7 -24 21 -16
4 U26A
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 24 0
1 U
8585 0 0
2
5.8987e-315 0
0
5 4071~
219 1729 647 0 3 22
0 12 11 13
0
0 0 624 90
4 4071
-7 -24 21 -16
4 U30A
25 -3 53 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 25 0
1 U
8809 0 0
2
43429.4 2
0
5 4081~
219 320 1137 0 3 22
0 17 16 14
0
0 0 624 512
4 4081
-7 -24 21 -16
4 U24A
-16 -25 12 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 21 0
1 U
5993 0 0
2
5.8987e-315 5.44228e-315
0
5 4073~
219 404 1195 0 4 22
0 5 4 3 16
0
0 0 624 512
4 4073
-7 -24 21 -16
4 U14B
-16 -25 12 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
8654 0 0
2
5.8987e-315 5.44487e-315
0
5 4082~
219 405 1091 0 5 22
0 10 9 8 6 17
0
0 0 624 512
4 4082
-7 -24 21 -16
4 U22A
-16 -28 12 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
7223 0 0
2
5.8987e-315 5.44746e-315
0
14 Logic Display~
6 1934 534 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
5.8987e-315 5.45005e-315
0
5 4081~
219 1681 870 0 3 22
0 21 20 19
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U18A
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
3104 0 0
2
5.8987e-315 5.45264e-315
0
5 4081~
219 1937 963 0 3 22
0 22 20 18
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U17A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 13 0
1 U
3296 0 0
2
5.8987e-315 5.45523e-315
0
14 Logic Display~
6 1641 1282 0 1 2
12 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
5.8987e-315 5.45782e-315
0
5 4049~
219 1621 1298 0 2 22
0 20 11
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 12 0
1 U
949 0 0
2
5.8987e-315 5.46041e-315
0
5 4081~
219 1531 549 0 3 22
0 33 9 32
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 18 0
1 U
3371 0 0
2
5.8987e-315 5.463e-315
0
5 4027~
219 1584 714 0 7 32
0 15 32 31 32 14 73 10
0
0 0 4720 0
4 4027
7 -60 35 -52
4 U27B
19 -61 47 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 23 0
1 U
7311 0 0
2
5.8987e-315 5.46559e-315
0
4 4585
219 849 1589 0 14 29
0 10 9 7 6 30 29 28 27 26
39 26 37 40 35
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U29
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 0 1 0 0 0
1 U
3409 0 0
2
5.8987e-315 5.46818e-315
0
4 4585
219 1474 1599 0 14 29
0 5 4 2 26 25 24 23 26 35
40 37 38 74 75
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U28
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
3526 0 0
2
5.8987e-315 5.47077e-315
0
5 4069~
219 877 1690 0 2 22
0 26 39
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
4129 0 0
2
5.8987e-315 5.47207e-315
0
5 4071~
219 1558 1655 0 3 22
0 38 37 36
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
6278 0 0
2
5.8987e-315 5.47336e-315
0
5 4081~
219 1609 1612 0 3 22
0 36 34 20
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U19C
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 18 0
1 U
3482 0 0
2
5.8987e-315 5.47466e-315
0
5 4049~
219 1631 1659 0 2 22
0 35 34
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U25F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 22 0
1 U
8323 0 0
2
5.8987e-315 5.47595e-315
0
14 Logic Display~
6 1732 532 0 1 2
12 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
43429.4 3
0
5 4049~
219 1737 797 0 2 22
0 18 42
0
0 0 624 602
4 4049
-7 -24 21 -16
4 U13A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 17 0
1 U
7622 0 0
2
43429.4 4
0
5 4049~
219 1719 796 0 2 22
0 21 43
0
0 0 624 602
4 4049
-7 -24 21 -16
4 U23F
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 19 0
1 U
816 0 0
2
43429.4 5
0
5 4081~
219 1732 755 0 3 22
0 43 42 12
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U21C
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 16 0
1 U
4656 0 0
2
43429.4 6
0
5 4081~
219 1610 838 0 3 22
0 45 46 21
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U21B
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 16 0
1 U
6356 0 0
2
5.8987e-315 5.47854e-315
0
14 Logic Display~
6 1833 527 0 1 2
11 19
0
0 0 53872 512
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7479 0 0
2
5.8987e-315 5.47984e-315
0
5 4049~
219 519 879 0 2 22
0 48 47
0
0 0 624 512
4 4049
-7 -24 21 -16
4 U15A
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
5690 0 0
2
43429.4 7
0
9 8-In NOR~
219 580 879 0 9 19
0 15 10 2 4 5 6 7 9 48
0
0 0 624 512
4 4078
-7 -24 21 -16
3 U12
3 -44 24 -36
0
15 DVDD=14;DGND=7;
97 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 2 3 4 5 9 10 11 12 13
2 3 4 5 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
5617 0 0
2
43429.4 8
0
5 4071~
219 386 741 0 3 22
0 49 47 45
0
0 0 624 90
4 4071
-7 -24 21 -16
3 U9B
28 -3 49 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
3903 0 0
2
43429.4 9
0
14 Logic Display~
6 1925 841 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4452 0 0
2
5.8987e-315 5.48113e-315
0
5 4049~
219 1632 1066 0 2 22
0 46 50
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
6282 0 0
2
5.8987e-315 5.48243e-315
0
5 4049~
219 1641 1216 0 2 22
0 53 52
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
7187 0 0
2
5.8987e-315 5.48372e-315
0
5 4081~
219 1619 1169 0 3 22
0 54 52 46
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U10A
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
6866 0 0
2
5.8987e-315 5.48502e-315
0
5 4071~
219 1568 1212 0 3 22
0 56 55 54
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
7670 0 0
2
5.8987e-315 5.48631e-315
0
14 Logic Display~
6 1547 1074 0 1 2
10 57
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
951 0 0
2
5.8987e-315 5.48761e-315
0
5 4069~
219 887 1247 0 2 22
0 59 58
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 6 0
1 U
9536 0 0
2
5.8987e-315 5.4889e-315
0
4 4585
219 1484 1156 0 14 29
0 4 2 59 59 62 61 59 59 53
60 55 56 76 57
0
0 0 4848 0
4 4585
-14 -60 14 -52
2 U7
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
5495 0 0
2
5.8987e-315 5.4902e-315
0
4 4585
219 859 1146 0 14 29
0 9 7 6 5 63 64 65 44 59
58 59 55 60 53
0
0 0 4848 0
4 4585
-14 -60 14 -52
2 U6
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 0 1 0 0 0
1 U
8152 0 0
2
5.8987e-315 5.49149e-315
0
5 4049~
219 1250 973 0 2 22
0 5 77
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5D
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 4 5 0
1 U
6223 0 0
2
5.8987e-315 5.49279e-315
0
5 4049~
219 1112 962 0 2 22
0 6 78
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5C
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 3 5 0
1 U
5441 0 0
2
5.8987e-315 5.49408e-315
0
5 4049~
219 962 957 0 2 22
0 7 79
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5B
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 2 5 0
1 U
3189 0 0
2
5.8987e-315 5.49538e-315
0
5 4049~
219 772 950 0 2 22
0 9 80
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5A
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 1 5 0
1 U
8460 0 0
2
5.8987e-315 5.49667e-315
0
14 Logic Display~
6 1480 984 0 1 2
10 2
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5179 0 0
2
5.8987e-315 5.49797e-315
0
14 Logic Display~
6 1414 986 0 1 2
10 4
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3593 0 0
2
5.8987e-315 5.49926e-315
0
14 Logic Display~
6 1296 987 0 1 2
10 5
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3928 0 0
2
5.8987e-315 5.50056e-315
0
14 Logic Display~
6 1178 988 0 1 2
10 6
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
363 0 0
2
5.8987e-315 5.50185e-315
0
14 Logic Display~
6 1039 983 0 1 2
10 7
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8132 0 0
2
5.8987e-315 5.50315e-315
0
14 Logic Display~
6 843 984 0 1 2
10 9
0
0 0 53872 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
65 0 0
2
5.8987e-315 5.50444e-315
0
5 4081~
219 1397 545 0 3 22
0 66 7 33
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
6609 0 0
2
5.8987e-315 5.50574e-315
0
5 4081~
219 1301 546 0 3 22
0 67 6 66
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
8995 0 0
2
5.8987e-315 5.50703e-315
0
5 4027~
219 1462 709 0 7 32
0 15 33 31 33 14 81 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U4B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 4 0
1 U
3918 0 0
2
5.8987e-315 5.50833e-315
0
5 4027~
219 1356 711 0 7 32
0 15 66 31 66 14 82 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U4A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
7519 0 0
2
5.8987e-315 5.50963e-315
0
5 4081~
219 1166 544 0 3 22
0 69 5 67
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
377 0 0
2
5.8987e-315 5.51092e-315
0
5 4081~
219 1039 552 0 3 22
0 2 4 69
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
8816 0 0
2
5.8987e-315 5.51222e-315
0
14 Logic Display~
6 808 493 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3877 0 0
2
5.8987e-315 5.51286e-315
0
5 4027~
219 1122 709 0 7 32
0 15 69 31 69 14 83 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
926 0 0
2
5.8987e-315 5.51351e-315
0
5 4027~
219 1256 711 0 7 32
0 15 67 31 67 14 84 6
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7262 0 0
2
5.8987e-315 5.51416e-315
0
5 4027~
219 988 718 0 7 32
0 15 2 31 2 14 85 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
5267 0 0
2
5.8987e-315 5.51481e-315
0
5 4027~
219 854 716 0 7 32
0 15 68 31 68 14 86 2
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
8838 0 0
2
5.8987e-315 5.51545e-315
0
5 4049~
219 1395 937 0 2 22
0 4 87
0
0 0 624 512
4 4049
-7 -24 21 -16
4 U11A
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 1 9 0
1 U
7159 0 0
2
5.8987e-315 5.5161e-315
0
5 4049~
219 1461 917 0 2 22
0 2 88
0
0 0 624 512
4 4049
-7 -24 21 -16
4 U11B
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 2 9 0
1 U
5812 0 0
2
5.8987e-315 5.51675e-315
0
5 4073~
219 524 487 0 4 22
0 51 41 45 31
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
331 0 0
2
5.8987e-315 5.5174e-315
0
5 4081~
219 1859 942 0 3 22
0 50 45 22
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U20D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 15 0
1 U
9604 0 0
2
5.8987e-315 5.51804e-315
0
173
0 1 2 0 0 12288 0 0 21 113 0 6
1452 1064
1287 1064
1287 1398
483 1398
483 1204
458 1204
2 3 3 0 0 4224 0 21 25 0 0 2
422 1204
424 1204
0 2 4 0 0 12288 0 0 25 126 0 6
1360 1047
1318 1047
1318 1378
516 1378
516 1195
424 1195
0 1 5 0 0 4096 0 0 25 118 0 4
803 1071
507 1071
507 1186
424 1186
0 4 6 0 0 4096 0 0 26 119 0 4
810 1047
494 1047
494 1105
425 1105
0 1 7 0 0 4096 0 0 22 120 0 6
996 1000
697 1000
697 1038
471 1038
471 1096
458 1096
2 3 8 0 0 4224 0 22 26 0 0 2
422 1096
425 1096
0 2 9 0 0 12288 0 0 26 121 0 6
823 993
671 993
671 1023
440 1023
440 1087
425 1087
0 1 10 0 0 8192 0 0 26 39 0 4
648 857
648 1010
425 1010
425 1078
1 2 11 0 0 8320 0 30 23 0 0 3
1641 1300
1741 1300
1741 663
3 1 12 0 0 4224 0 43 23 0 0 3
1731 731
1731 663
1723 663
3 1 13 0 0 12416 0 23 40 0 0 4
1732 617
1732 619
1732 619
1732 550
3 5 14 0 0 8320 0 24 78 0 0 5
295 1137
295 816
820 816
820 722
854 722
1 0 15 0 0 4096 0 78 0 0 87 2
854 659
739 659
4 2 16 0 0 8320 0 25 24 0 0 3
379 1195
340 1195
340 1146
5 1 17 0 0 8320 0 26 24 0 0 4
380 1091
349 1091
349 1128
340 1128
0 1 18 0 0 8320 0 0 27 21 0 3
1939 859
1934 859
1934 552
3 1 19 0 0 8320 0 28 45 0 0 3
1680 846
1833 846
1833 545
0 2 20 0 0 4096 0 0 28 22 0 3
1913 1041
1689 1041
1689 891
0 1 21 0 0 4096 0 0 28 65 0 3
1653 814
1653 891
1671 891
3 1 18 0 0 0 0 29 49 0 0 3
1958 963
1958 859
1925 859
0 2 20 0 0 8320 0 0 29 50 0 3
1608 1350
1913 1350
1913 972
3 1 22 0 0 4224 0 82 29 0 0 3
1880 942
1913 942
1913 954
1 2 11 0 0 0 0 30 31 0 0 3
1641 1300
1641 1298
1642 1298
0 3 2 0 0 0 0 0 35 131 0 4
1480 952
1345 952
1345 1581
1442 1581
0 1 5 0 0 8192 0 0 35 133 0 4
1296 948
1232 948
1232 1563
1442 1563
0 4 6 0 0 12416 0 0 34 128 0 7
1157 962
1157 940
582 940
582 1520
768 1520
768 1580
817 1580
0 3 7 0 0 12416 0 0 34 129 0 7
1010 957
1010 930
607 930
607 1503
788 1503
788 1571
817 1571
0 2 9 0 0 12288 0 0 34 130 0 7
807 950
807 923
625 923
625 1488
805 1488
805 1562
817 1562
0 1 10 0 0 12416 0 0 34 39 0 5
1644 682
2043 682
2043 1500
817 1500
817 1553
1 7 23 0 0 4224 0 1 35 0 0 4
653 1798
1392 1798
1392 1617
1442 1617
1 6 24 0 0 4224 0 6 35 0 0 4
653 1766
1372 1766
1372 1608
1442 1608
1 5 25 0 0 4224 0 5 35 0 0 4
655 1728
1349 1728
1349 1599
1442 1599
0 0 26 0 0 4096 0 0 0 61 62 2
1418 1602
1418 1630
1 8 27 0 0 12416 0 8 34 0 0 4
659 1689
734 1689
734 1616
817 1616
1 7 28 0 0 12416 0 2 34 0 0 4
659 1642
672 1642
672 1607
817 1607
1 6 29 0 0 4224 0 3 34 0 0 4
662 1585
743 1585
743 1598
817 1598
1 5 30 0 0 4224 0 4 34 0 0 4
661 1538
757 1538
757 1589
817 1589
7 2 10 0 0 0 0 33 47 0 0 6
1608 678
1644 678
1644 768
1454 768
1454 857
609 857
0 3 31 0 0 4096 0 0 33 141 0 4
1408 592
1534 592
1534 687
1560 687
2 4 32 0 0 8192 0 33 33 0 0 4
1560 678
1546 678
1546 696
1560 696
3 2 32 0 0 8320 0 32 33 0 0 3
1552 549
1560 549
1560 678
0 2 9 0 0 0 0 0 32 136 0 3
1508 673
1507 673
1507 558
0 1 33 0 0 4096 0 0 32 138 0 3
1429 545
1507 545
1507 540
1 1 15 0 0 4096 0 70 33 0 0 3
1462 652
1584 652
1584 657
5 5 14 0 0 0 0 70 33 0 0 3
1462 715
1462 720
1584 720
0 2 4 0 0 0 0 0 35 126 0 3
1386 1003
1386 1572
1442 1572
2 2 34 0 0 8320 0 39 38 0 0 3
1652 1659
1652 1633
1617 1633
0 1 35 0 0 8192 0 0 39 60 0 5
1436 1644
1436 1633
1605 1633
1605 1659
1616 1659
1 3 20 0 0 0 0 31 38 0 0 3
1606 1298
1608 1298
1608 1588
1 3 36 0 0 4224 0 38 37 0 0 3
1599 1633
1599 1655
1591 1655
0 2 37 0 0 8192 0 0 37 58 0 4
1438 1662
1438 1683
1545 1683
1545 1664
12 1 38 0 0 4224 0 35 37 0 0 3
1506 1617
1545 1617
1545 1646
2 10 39 0 0 8320 0 36 34 0 0 3
898 1690
898 1643
817 1643
0 1 26 0 0 0 0 0 36 57 0 3
849 1689
849 1690
862 1690
0 9 26 0 0 8192 0 0 34 57 0 4
817 1663
791 1663
791 1634
817 1634
0 11 26 0 0 4096 0 0 34 62 0 4
849 1707
849 1672
817 1672
817 1652
12 11 37 0 0 12416 0 34 35 0 0 4
881 1607
1160 1607
1160 1662
1442 1662
13 10 40 0 0 4224 0 34 35 0 0 4
881 1598
1180 1598
1180 1653
1442 1653
14 9 35 0 0 4224 0 34 35 0 0 4
881 1589
1191 1589
1191 1644
1442 1644
0 4 26 0 0 0 0 0 35 0 0 3
1418 1610
1418 1590
1442 1590
1 8 26 0 0 4224 0 7 35 0 0 4
832 1707
1418 1707
1418 1626
1442 1626
1 2 41 0 0 4224 0 10 81 0 0 4
333 471
492 471
492 487
500 487
1 1 18 0 0 0 0 49 41 0 0 3
1925 859
1740 859
1740 815
3 1 21 0 0 4224 0 44 42 0 0 2
1609 814
1722 814
2 2 42 0 0 4224 0 41 43 0 0 4
1740 779
1740 770
1740 770
1740 776
2 1 43 0 0 12416 0 42 43 0 0 4
1722 778
1722 779
1722 779
1722 776
1 0 44 0 0 0 0 9 0 0 125 2
669 1246
669 1246
0 2 45 0 0 8192 0 0 82 70 0 3
1566 859
1566 951
1835 951
0 1 45 0 0 12416 0 0 44 81 0 6
389 675
518 675
518 839
1538 839
1538 859
1600 859
2 0 46 0 0 0 0 44 0 0 99 2
1618 859
1618 859
2 2 47 0 0 8320 0 46 48 0 0 3
504 879
398 879
398 757
9 1 48 0 0 4224 0 47 46 0 0 2
553 879
540 879
8 0 9 0 0 0 0 47 0 0 93 2
609 911
609 911
7 0 7 0 0 0 0 47 0 0 92 2
609 902
609 902
6 0 6 0 0 0 0 47 0 0 91 2
609 893
609 893
5 0 5 0 0 0 0 47 0 0 90 2
609 884
609 884
4 0 4 0 0 0 0 47 0 0 89 2
609 875
609 875
3 0 2 0 0 0 0 47 0 0 88 2
609 866
609 866
1 0 15 0 0 0 0 47 0 0 87 2
609 848
609 848
3 3 45 0 0 0 0 48 81 0 0 3
389 711
389 496
500 496
1 1 49 0 0 20608 0 11 48 0 0 6
166 971
231 971
231 881
230 881
230 757
380 757
2 1 50 0 0 8320 0 50 82 0 0 4
1653 1066
1718 1066
1718 933
1835 933
4 0 31 0 0 4224 0 81 0 0 86 4
545 487
781 487
781 522
808 522
3 1 51 0 0 12416 0 20 81 0 0 5
336 409
409 409
409 425
500 425
500 478
1 0 31 0 0 0 0 74 0 0 152 2
808 511
808 524
1 0 15 0 0 4224 0 19 0 0 0 3
739 651
739 848
603 848
0 0 2 0 0 4224 0 0 0 0 131 2
603 866
1481 866
0 0 4 0 0 4224 0 0 0 0 132 2
603 875
1415 875
0 0 5 0 0 4224 0 0 0 0 133 2
603 884
1298 884
0 0 6 0 0 0 0 0 0 0 134 2
603 893
1171 893
0 0 7 0 0 0 0 0 0 0 135 2
603 902
1038 902
0 0 9 0 0 0 0 0 0 0 136 2
603 911
882 911
1 0 2 0 0 0 0 80 0 0 131 2
1482 917
1481 917
1 0 4 0 0 0 0 79 0 0 132 2
1416 937
1415 937
1 0 46 0 0 4096 0 50 0 0 99 2
1617 1066
1618 1066
2 2 52 0 0 8320 0 51 52 0 0 3
1662 1216
1662 1190
1627 1190
0 1 53 0 0 8192 0 0 51 110 0 5
1446 1201
1446 1190
1615 1190
1615 1216
1626 1216
0 3 46 0 0 4224 0 0 52 0 0 2
1618 854
1618 1145
1 3 54 0 0 4224 0 52 53 0 0 3
1609 1190
1609 1212
1601 1212
0 2 55 0 0 8192 0 0 53 108 0 4
1448 1219
1448 1240
1555 1240
1555 1221
12 1 56 0 0 4224 0 56 53 0 0 3
1516 1174
1555 1174
1555 1203
14 1 57 0 0 8320 0 56 54 0 0 3
1516 1156
1547 1156
1547 1092
2 10 58 0 0 8320 0 55 57 0 0 3
908 1247
908 1200
827 1200
0 1 59 0 0 8192 0 0 55 107 0 3
859 1246
859 1247
872 1247
0 9 59 0 0 8192 0 0 57 107 0 4
827 1220
801 1220
801 1191
827 1191
0 11 59 0 0 4096 0 0 57 117 0 4
859 1264
859 1229
827 1229
827 1209
12 11 55 0 0 12416 0 57 56 0 0 4
891 1164
1170 1164
1170 1219
1452 1219
13 10 60 0 0 4224 0 57 56 0 0 4
891 1155
1190 1155
1190 1210
1452 1210
14 9 53 0 0 4224 0 57 56 0 0 4
891 1146
1201 1146
1201 1201
1452 1201
1 6 61 0 0 4224 0 13 56 0 0 4
663 1323
1434 1323
1434 1165
1452 1165
1 5 62 0 0 4224 0 14 56 0 0 4
665 1285
1440 1285
1440 1156
1452 1156
0 2 2 0 0 0 0 0 56 131 0 3
1480 964
1452 964
1452 1129
0 3 59 0 0 0 0 0 56 115 0 3
1428 1147
1428 1138
1452 1138
0 4 59 0 0 0 0 0 56 116 0 3
1428 1174
1428 1147
1452 1147
0 7 59 0 0 0 0 0 56 117 0 3
1428 1183
1428 1174
1452 1174
1 8 59 0 0 4224 0 12 56 0 0 4
842 1264
1428 1264
1428 1183
1452 1183
0 4 5 0 0 0 0 0 57 127 0 5
1281 973
1281 1058
803 1058
803 1137
827 1137
0 3 6 0 0 0 0 0 57 128 0 5
1149 962
1149 1034
810 1034
810 1128
827 1128
0 2 7 0 0 0 0 0 57 129 0 5
996 957
996 1022
817 1022
817 1119
827 1119
0 1 9 0 0 0 0 0 57 130 0 3
823 950
823 1110
827 1110
1 5 63 0 0 4224 0 15 57 0 0 4
671 1095
793 1095
793 1146
827 1146
1 6 64 0 0 4224 0 16 57 0 0 4
672 1142
777 1142
777 1155
827 1155
1 7 65 0 0 4224 0 17 57 0 0 4
669 1199
751 1199
751 1164
827 1164
0 8 44 0 0 4224 0 0 57 0 0 4
665 1246
761 1246
761 1173
827 1173
0 1 4 0 0 0 0 0 56 132 0 6
1414 956
1396 956
1396 1003
1360 1003
1360 1120
1452 1120
1 1 5 0 0 0 0 64 58 0 0 2
1296 973
1271 973
0 1 6 0 0 0 0 0 59 134 0 3
1178 961
1178 962
1133 962
0 1 7 0 0 0 0 0 60 135 0 2
1039 957
983 957
0 1 9 0 0 0 0 0 61 136 0 3
843 952
843 950
793 950
0 1 2 0 0 0 0 0 62 170 0 6
894 682
894 830
1481 830
1481 942
1480 942
1480 970
7 1 4 0 0 0 0 77 63 0 0 7
1012 682
1051 682
1051 785
1415 785
1415 946
1414 946
1414 972
7 1 5 0 0 0 0 75 64 0 0 7
1146 673
1162 673
1162 806
1298 806
1298 944
1296 944
1296 973
7 1 6 0 0 0 0 76 65 0 0 6
1280 675
1280 856
1171 856
1171 940
1178 940
1178 974
7 1 7 0 0 0 0 71 66 0 0 6
1380 675
1380 760
1038 760
1038 940
1039 940
1039 969
7 1 9 0 0 12416 0 70 67 0 0 7
1486 673
1517 673
1517 745
882 745
882 941
843 941
843 970
0 4 33 0 0 0 0 0 70 138 0 3
1431 672
1431 691
1438 691
3 2 33 0 0 8320 0 68 70 0 0 4
1418 545
1431 545
1431 673
1438 673
3 1 66 0 0 8192 0 69 68 0 0 3
1322 546
1322 536
1373 536
7 2 7 0 0 0 0 71 68 0 0 4
1380 675
1380 567
1373 567
1373 554
0 3 31 0 0 0 0 0 70 146 0 4
1298 592
1409 592
1409 682
1438 682
5 5 14 0 0 0 0 71 70 0 0 3
1356 717
1356 715
1462 715
1 1 15 0 0 0 0 71 70 0 0 3
1356 654
1356 652
1462 652
5 5 14 0 0 0 0 76 71 0 0 2
1256 717
1356 717
1 1 15 0 0 0 0 76 71 0 0 2
1256 654
1356 654
0 3 31 0 0 0 0 0 71 171 0 4
1212 592
1298 592
1298 684
1332 684
0 4 66 0 0 0 0 0 71 148 0 3
1322 675
1322 693
1332 693
3 2 66 0 0 4224 0 69 71 0 0 3
1322 546
1322 675
1332 675
3 1 67 0 0 8192 0 72 69 0 0 3
1187 544
1187 537
1277 537
7 2 6 0 0 0 0 76 69 0 0 3
1280 675
1277 675
1277 555
0 3 31 0 0 0 0 0 78 173 0 3
815 592
815 689
830 689
0 0 31 0 0 0 0 0 0 0 173 2
808 515
808 592
0 4 68 0 0 8192 0 0 78 154 0 3
754 680
754 698
830 698
1 2 68 0 0 8320 0 18 78 0 0 4
749 584
754 584
754 680
830 680
5 5 14 0 0 0 0 75 76 0 0 3
1122 715
1122 717
1256 717
5 5 14 0 0 0 0 77 75 0 0 3
988 724
1122 724
1122 715
5 5 14 0 0 0 0 78 77 0 0 3
854 722
854 724
988 724
1 1 15 0 0 0 0 75 76 0 0 3
1122 652
1122 654
1256 654
1 1 15 0 0 0 0 77 75 0 0 4
988 661
1101 661
1101 652
1122 652
1 1 15 0 0 0 0 78 77 0 0 3
854 659
854 661
988 661
0 4 67 0 0 0 0 0 76 162 0 3
1187 675
1187 693
1232 693
3 2 67 0 0 4224 0 72 76 0 0 3
1187 544
1187 675
1232 675
3 1 69 0 0 8192 0 73 72 0 0 3
1060 552
1060 535
1142 535
7 2 5 0 0 0 0 75 72 0 0 3
1146 673
1142 673
1142 553
0 4 69 0 0 0 0 0 75 166 0 3
1060 672
1060 691
1098 691
3 2 69 0 0 4224 0 73 75 0 0 3
1060 552
1060 673
1098 673
7 2 4 0 0 0 0 77 73 0 0 3
1012 682
1015 682
1015 561
0 1 2 0 0 0 0 0 73 170 0 3
906 682
906 543
1015 543
0 4 2 0 0 0 0 0 77 170 0 3
926 682
926 700
964 700
7 2 2 0 0 0 0 78 77 0 0 3
878 680
878 682
964 682
0 3 31 0 0 0 0 0 76 172 0 4
1073 592
1212 592
1212 684
1232 684
0 3 31 0 0 0 0 0 75 173 0 4
944 592
1073 592
1073 682
1098 682
0 3 31 0 0 0 0 0 77 0 0 4
802 592
946 592
946 691
964 691
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1680 1296 1827 1320
1685 1298 1821 1314
17 pelo tempo m�nimo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 42
1680 1279 2027 1303
1685 1281 2021 1297
42 Controle interno que mostra o sinal aberto
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
1769 459 1887 478
1781 464 1874 477
14 Luzes do sinal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
52 993 263 1017
57 995 257 1011
25 Input para fechar o sinal
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
665 643 698 667
669 645 693 661
3 GND
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
668 572 703 596
673 574 697 590
3 VCC
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
