CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 40 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
66
13 Logic Switch~
5 89 1860 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V23
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8628 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 88 1922 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3516 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 86 1708 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7639 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 97 1488 0 1 11
0 23
0
0 0 21344 0
2 0V
-1 -13 13 -5
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
468 0 0
2
5.89862e-315 5.32571e-315
0
13 Logic Switch~
5 96 1537 0 1 11
0 21
0
0 0 21344 0
2 0V
-1 -13 13 -5
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
360 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 88 1597 0 1 11
0 20
0
0 0 21344 0
2 0V
-1 -13 13 -5
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7326 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 87 1646 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3479 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 102 1284 0 1 11
0 30
0
0 0 21344 0
2 0V
-1 -13 13 -5
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7329 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 107 1233 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3530 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 101 1333 0 1 11
0 32
0
0 0 21344 0
2 0V
-1 -13 13 -5
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8542 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 138 1116 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3445 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 155 1025 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V12
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9600 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 160 958 0 10 11
0 38 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5719 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 145 843 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3686 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 159 563 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
861 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 154 630 0 10 11
0 45 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5536 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 153 678 0 10 11
0 44 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6385 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 178 443 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9434 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 179 395 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8462 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 184 328 0 10 11
0 55 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-1 -13 13 -5
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3388 0 0
2
5.89862e-315 0
0
13 Logic Switch~
5 185 194 0 10 11
0 59 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-10 -14 4 -6
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
7552 0 0
2
5.89862e-315 5.26354e-315
0
13 Logic Switch~
5 183 141 0 1 11
0 57
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3634 0 0
2
5.89862e-315 5.30499e-315
0
13 Logic Switch~
5 189 91 0 1 11
0 58
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4841 0 0
2
5.89862e-315 5.32571e-315
0
8 Battery~
219 490 1808 0 2 5
0 3 60
0
0 0 864 180
2 5V
13 0 27 8
3 V24
11 -12 32 -4
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 512 1 0 0 0
1 V
7680 0 0
2
5.89862e-315 0
0
4 LED~
171 488 1857 0 2 2
10 3 4
0
0 0 880 0
4 LED0
17 0 45 8
2 D4
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3220 0 0
2
5.89862e-315 0
0
5 4001~
219 393 1849 0 3 22
0 8 5 4
0
0 0 608 0
4 4001
-14 -24 14 -16
3 U6C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 12 0
1 U
3230 0 0
2
5.89862e-315 0
0
5 4081~
219 306 1920 0 3 22
0 10 9 5
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 19 0
1 U
7598 0 0
2
5.89862e-315 0
0
5 4049~
219 264 1930 0 2 22
0 6 9
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U7D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 17 0
1 U
7184 0 0
2
5.89862e-315 0
0
5 4049~
219 263 1911 0 2 22
0 7 10
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 17 0
1 U
5144 0 0
2
5.89862e-315 0
0
5 4081~
219 239 1835 0 3 22
0 7 6 8
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 19 0
1 U
6284 0 0
2
5.89862e-315 0
0
9 Inverter~
13 519 1509 0 2 22
0 11 16
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U13D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 23 0
1 U
3779 0 0
2
5.89862e-315 0
0
9 Inverter~
13 520 1500 0 2 22
0 13 17
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U13C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 23 0
1 U
9382 0 0
2
5.89862e-315 0
0
9 Inverter~
13 519 1491 0 2 22
0 14 18
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U13B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 23 0
1 U
5951 0 0
2
5.89862e-315 0
0
9 Inverter~
13 521 1482 0 2 22
0 15 19
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U13A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 23 0
1 U
9697 0 0
2
5.89862e-315 0
0
8 4-In OR~
219 555 1495 0 5 22
0 19 18 17 16 61
0
0 0 608 0
4 4072
-14 -24 14 -16
4 U12A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 22 0
1 U
3832 0 0
2
5.89862e-315 0
0
9 Inverter~
13 285 1696 0 2 22
0 12 11
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U11F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 21 0
1 U
3648 0 0
2
5.89862e-315 0
0
9 Inverter~
13 192 1437 0 2 22
0 23 22
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U11E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 21 0
1 U
3124 0 0
2
5.89862e-315 0
0
9 Inverter~
13 285 1541 0 2 22
0 20 24
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U11D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 21 0
1 U
834 0 0
2
5.89862e-315 0
0
9 Inverter~
13 283 1524 0 2 22
0 21 25
0
0 0 608 0
5 74F04
-18 -19 17 -11
4 U11C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 21 0
1 U
6448 0 0
2
5.89862e-315 0
0
5 4011~
219 326 1532 0 3 22
0 25 24 14
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 20 0
1 U
6517 0 0
2
5.89862e-315 0
0
5 4011~
219 338 1437 0 3 22
0 22 21 15
0
0 0 608 0
4 4011
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 20 0
1 U
7298 0 0
2
5.89862e-315 0
0
4 LED~
171 356 1286 0 2 2
10 26 27
0
0 0 880 0
4 LED0
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
9836 0 0
2
5.89862e-315 0
0
5 4049~
219 166 1333 0 2 22
0 32 31
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U7B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 17 0
1 U
3111 0 0
2
5.89862e-315 0
0
5 4071~
219 208 1319 0 3 22
0 30 31 29
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
6852 0 0
2
5.89862e-315 0
0
5 4081~
219 224 1244 0 3 22
0 28 29 26
0
0 0 608 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 19 0
1 U
5866 0 0
2
5.89862e-315 0
0
10 2-In NAND~
219 523 1018 0 3 22
0 35 33 62
0
0 0 608 0
5 74F37
-10 -24 25 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 18 0
1 U
3461 0 0
2
5.89862e-315 0
0
5 4001~
219 380 1082 0 3 22
0 34 36 33
0
0 0 608 0
4 4001
-14 -24 14 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 12 0
1 U
4744 0 0
2
5.89862e-315 0
0
5 4049~
219 272 1115 0 2 22
0 37 36
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 17 0
1 U
7721 0 0
2
5.89862e-315 0
0
5 4001~
219 316 989 0 3 22
0 38 34 35
0
0 0 608 0
4 4001
-14 -24 14 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 12 0
1 U
368 0 0
2
5.89862e-315 0
0
9 3-In AND~
219 377 792 0 4 22
0 43 40 39 46
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 15 0
1 U
4982 0 0
2
5.89862e-315 0
0
9 3-In AND~
219 386 703 0 4 22
0 42 40 41 47
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 16 0
1 U
7855 0 0
2
5.89862e-315 0
0
8 3-In OR~
219 489 629 0 4 22
0 48 47 46 63
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 2 13 0
1 U
4170 0 0
2
5.89862e-315 0
0
9 3-In AND~
219 383 590 0 4 22
0 43 40 41 48
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 16 0
1 U
3791 0 0
2
5.89862e-315 0
0
5 4049~
219 272 680 0 2 22
0 44 41
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 11 0
1 U
331 0 0
2
5.89862e-315 0
0
5 4049~
219 272 571 0 2 22
0 42 43
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 11 0
1 U
8783 0 0
2
5.89862e-315 5.26354e-315
0
5 4049~
219 271 624 0 2 22
0 45 40
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
9888 0 0
2
5.89862e-315 0
0
7 Ground~
168 604 389 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6667 0 0
2
5.89862e-315 0
0
4 LED~
171 604 374 0 2 2
10 2 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8701 0 0
2
5.89862e-315 0
0
9 3-In AND~
219 584 365 0 4 22
0 51 50 49 2
0
0 0 608 0
5 74F11
-18 -28 17 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 16 0
1 U
7651 0 0
2
5.89862e-315 0
0
5 4071~
219 397 321 0 3 22
0 54 53 52
0
0 0 608 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
5986 0 0
2
5.89862e-315 0
0
5 4049~
219 482 319 0 2 22
0 52 51
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
4267 0 0
2
5.89862e-315 0
0
5 4049~
219 319 351 0 2 22
0 50 53
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
7787 0 0
2
5.89862e-315 0
0
5 4049~
219 320 298 0 2 22
0 55 54
0
0 0 608 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
4802 0 0
2
5.89862e-315 0
0
8 3-In OR~
219 364 141 0 4 22
0 58 57 56 2
0
0 0 608 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
7867 0 0
2
5.89862e-315 0
0
7 Ground~
168 566 128 0 1 3
0 2
0
0 0 53344 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3797 0 0
2
43359.9 0
0
4 LED~
171 566 147 0 2 2
10 2 2
0
0 0 880 0
4 LED0
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7294 0 0
2
43359.9 1
0
74
1 1 3 0 0 4224 0 25 24 0 0 2
488 1847
488 1817
3 2 4 0 0 4224 0 26 25 0 0 4
432 1849
460 1849
460 1867
488 1867
3 2 5 0 0 8320 0 27 26 0 0 3
327 1920
380 1920
380 1858
0 1 6 0 0 8192 0 0 28 6 0 3
187 1922
187 1930
249 1930
0 1 7 0 0 4224 0 0 29 8 0 3
180 1826
180 1911
248 1911
1 2 6 0 0 4224 0 2 30 0 0 4
100 1922
200 1922
200 1844
215 1844
3 1 8 0 0 4224 0 30 26 0 0 3
260 1835
380 1835
380 1840
1 1 7 0 0 0 0 1 30 0 0 4
101 1860
154 1860
154 1826
215 1826
2 2 9 0 0 8320 0 28 27 0 0 3
285 1930
285 1929
282 1929
2 1 10 0 0 4224 0 29 27 0 0 2
284 1911
282 1911
2 1 11 0 0 4224 0 36 31 0 0 3
306 1696
504 1696
504 1509
1 1 12 0 0 4224 0 36 3 0 0 3
270 1696
98 1696
98 1708
1 1 13 0 0 4224 0 7 32 0 0 4
99 1646
492 1646
492 1500
505 1500
3 1 14 0 0 4224 0 40 33 0 0 4
353 1532
486 1532
486 1491
504 1491
3 1 15 0 0 4224 0 41 34 0 0 3
365 1437
506 1437
506 1482
2 4 16 0 0 4224 0 31 35 0 0 2
540 1509
538 1509
2 3 17 0 0 4224 0 32 35 0 0 2
541 1500
538 1500
2 2 18 0 0 4224 0 33 35 0 0 2
540 1491
538 1491
2 1 19 0 0 4224 0 34 35 0 0 2
542 1482
538 1482
1 1 20 0 0 4224 0 6 38 0 0 3
100 1597
270 1597
270 1541
0 1 21 0 0 8192 0 0 39 22 0 3
147 1523
147 1524
268 1524
1 2 21 0 0 12416 0 5 41 0 0 4
108 1537
147 1537
147 1446
314 1446
2 1 22 0 0 4224 0 37 41 0 0 4
213 1437
304 1437
304 1428
314 1428
1 1 23 0 0 12416 0 4 37 0 0 4
109 1488
115 1488
115 1437
177 1437
2 2 24 0 0 4224 0 38 40 0 0 2
306 1541
302 1541
2 1 25 0 0 8320 0 39 40 0 0 3
304 1524
304 1523
302 1523
2 0 21 0 0 0 0 41 0 0 0 2
314 1446
320 1446
3 1 26 0 0 4224 0 45 42 0 0 3
245 1244
356 1244
356 1276
0 2 27 0 0 4224 0 0 42 0 0 2
356 1276
356 1296
1 1 28 0 0 8320 0 9 45 0 0 3
119 1233
119 1235
200 1235
3 2 29 0 0 4224 0 44 45 0 0 4
241 1319
241 1267
200 1267
200 1253
1 1 30 0 0 4224 0 8 44 0 0 3
114 1284
195 1284
195 1310
2 2 31 0 0 4224 0 43 44 0 0 3
187 1333
195 1333
195 1328
1 1 32 0 0 4224 0 10 43 0 0 2
113 1333
151 1333
3 2 33 0 0 4224 0 47 46 0 0 3
419 1082
499 1082
499 1027
0 1 34 0 0 8320 0 0 47 40 0 3
246 1025
246 1073
367 1073
3 1 35 0 0 4224 0 49 46 0 0 3
355 989
499 989
499 1009
2 2 36 0 0 4224 0 48 47 0 0 3
293 1115
367 1115
367 1091
1 1 37 0 0 8320 0 11 48 0 0 3
150 1116
150 1115
257 1115
1 2 34 0 0 0 0 12 49 0 0 4
167 1025
257 1025
257 998
303 998
1 1 38 0 0 4224 0 13 49 0 0 4
172 958
258 958
258 980
303 980
1 3 39 0 0 4224 0 14 50 0 0 3
157 843
353 843
353 801
0 2 40 0 0 4224 0 0 50 45 0 3
302 703
302 792
353 792
0 3 41 0 0 4096 0 0 51 48 0 3
332 680
332 712
362 712
0 2 40 0 0 0 0 0 51 50 0 3
302 624
302 703
362 703
0 1 42 0 0 8320 0 0 51 53 0 3
217 563
217 694
362 694
0 1 43 0 0 12416 0 0 50 52 0 5
312 571
312 512
97 512
97 783
353 783
2 3 41 0 0 8320 0 54 53 0 0 3
293 680
359 680
359 599
1 1 44 0 0 8320 0 17 54 0 0 3
165 678
165 680
257 680
2 2 40 0 0 0 0 56 53 0 0 4
292 624
347 624
347 590
359 590
1 1 45 0 0 4224 0 16 56 0 0 3
166 630
256 630
256 624
2 1 43 0 0 0 0 55 53 0 0 3
293 571
359 571
359 581
1 1 42 0 0 0 0 15 55 0 0 3
171 563
257 563
257 571
4 3 46 0 0 8320 0 50 52 0 0 3
398 792
476 792
476 638
4 2 47 0 0 4224 0 51 52 0 0 3
407 703
407 629
477 629
4 1 48 0 0 4224 0 53 52 0 0 3
404 590
476 590
476 620
1 0 2 0 0 0 0 57 0 0 59 2
604 383
604 383
1 4 2 0 0 4096 0 58 59 0 0 3
604 364
604 365
605 365
0 2 2 0 0 4096 0 0 58 58 0 2
604 364
604 384
1 3 49 0 0 4224 0 18 59 0 0 3
190 443
560 443
560 374
0 2 50 0 0 4224 0 0 59 64 0 4
304 377
466 377
466 365
560 365
2 1 51 0 0 4224 0 61 59 0 0 4
503 319
544 319
544 356
560 356
3 1 52 0 0 8320 0 60 61 0 0 3
430 321
430 319
467 319
1 1 50 0 0 0 0 19 62 0 0 3
191 395
304 395
304 351
2 2 53 0 0 4224 0 62 60 0 0 3
340 351
384 351
384 330
2 1 54 0 0 4224 0 63 60 0 0 3
341 298
384 298
384 312
1 1 55 0 0 4224 0 20 63 0 0 4
196 328
257 328
257 298
305 298
2 4 2 0 0 4224 0 66 64 0 0 4
566 157
453 157
453 141
397 141
0 3 56 0 0 4224 0 0 64 0 0 3
196 197
351 197
351 150
1 2 57 0 0 4224 0 22 64 0 0 5
195 141
332 141
332 142
352 142
352 141
1 1 58 0 0 4224 0 23 64 0 0 4
201 91
353 91
353 132
351 132
1 1 2 0 0 0 0 65 66 0 0 4
566 136
566 129
566 129
566 137
1 0 2 0 0 0 0 66 0 0 74 2
566 137
566 137
0 2 2 0 0 0 0 0 66 0 0 2
566 137
566 157
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
25 1745 130 1770
43 1753 111 1768
9 pagina 18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
43 27 123 66
49 29 116 59
9 Pagina 15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
30 911 110 950
36 913 103 943
9 Pagina 16
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
42 1163 120 1184
47 1166 114 1181
9 pagina 17
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
