CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 46 281 0 1 11
0 4
0
0 0 22384 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-26 -10 -19 -2
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6851 0 0
2
5.89797e-315 0
0
13 Logic Switch~
5 54 93 0 1 11
0 5
0
0 0 22384 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-22 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7156 0 0
2
5.89797e-315 0
0
4 LED~
171 434 209 0 2 2
10 3 2
0
0 0 864 90
4 LED1
-12 -21 16 -13
2 D2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8416 0 0
2
5.89797e-315 5.26354e-315
0
7 Ground~
168 455 207 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3383 0 0
2
5.89797e-315 0
0
10 2-In NAND~
219 365 211 0 3 22
0 8 7 3
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
398 0 0
2
5.89797e-315 0
0
10 2-In NAND~
219 287 274 0 3 22
0 6 4 7
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7742 0 0
2
5.89797e-315 0
0
10 2-In NAND~
219 225 64 0 3 22
0 5 6 8
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
5272 0 0
2
5.89797e-315 0
0
10 2-In NAND~
219 145 165 0 3 22
0 5 4 6
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
4993 0 0
2
5.89797e-315 0
0
10
2 1 2 0 0 12432 0 3 4 0 0 4
447 210
447 212
448 212
448 208
3 1 3 0 0 4224 0 5 3 0 0 4
392 211
411 211
411 210
427 210
0 2 4 0 0 8192 0 0 8 5 0 3
91 281
121 281
121 174
0 1 5 0 0 4096 0 0 8 10 0 3
122 55
122 156
121 156
1 2 4 0 0 12416 0 1 6 0 0 4
58 281
128 281
128 283
263 283
0 1 6 0 0 4224 0 0 6 7 0 3
200 113
200 265
263 265
2 3 6 0 0 128 0 7 8 0 0 6
201 73
202 73
202 113
200 113
200 165
172 165
3 2 7 0 0 8320 0 6 5 0 0 4
314 274
311 274
311 220
341 220
3 1 8 0 0 8320 0 7 5 0 0 4
252 64
311 64
311 202
341 202
1 1 5 0 0 12416 0 2 7 0 0 4
66 93
92 93
92 55
201 55
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
