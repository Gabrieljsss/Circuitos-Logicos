CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
176 86 1918 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 182 457 279
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 483 424 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43430.5 0
0
13 Logic Switch~
5 196 297 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43430.5 1
0
13 Logic Switch~
5 202 133 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43430.5 2
0
13 Logic Switch~
5 149 187 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -13 8 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.89871e-315 0
0
5 4049~
219 755 129 0 2 22
0 4 8
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5B
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
8157 0 0
2
43430.5 3
0
5 4081~
219 722 138 0 3 22
0 8 7 6
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
5572 0 0
2
43430.5 4
0
5 4071~
219 566 126 0 3 22
0 4 11 10
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
43430.5 5
0
5 4049~
219 324 300 0 2 22
0 7 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
7361 0 0
2
43430.5 6
0
5 4081~
219 492 107 0 3 22
0 3 11 13
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
4747 0 0
2
43430.5 7
0
5 4071~
219 348 96 0 3 22
0 2 13 12
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
972 0 0
2
43430.5 8
0
12 Hex Display~
7 956 230 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3472 0 0
2
43430.5 9
0
7 Pulser~
4 150 91 0 10 12
0 15 16 17 18 0 0 5 5 5
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9998 0 0
2
5.89871e-315 5.26354e-315
0
5 4027~
219 804 241 0 7 32
0 5 6 14 9 5 19 2
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3536 0 0
2
5.89871e-315 5.30499e-315
0
5 4027~
219 603 239 0 7 32
0 5 9 14 10 5 20 3
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4597 0 0
2
5.89871e-315 5.32571e-315
0
5 4027~
219 408 238 0 7 32
0 5 12 14 3 5 21 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3835 0 0
2
5.89871e-315 5.34643e-315
0
29
0 1 2 0 0 8192 0 0 11 16 0 5
828 198
901 198
901 293
965 293
965 254
0 2 3 0 0 4224 0 0 11 14 0 3
642 268
959 268
959 254
0 3 4 0 0 8320 0 0 11 5 0 6
432 124
432 33
927 33
927 264
953 264
953 254
0 1 4 0 0 0 0 0 5 5 0 4
531 121
531 41
776 41
776 129
7 1 4 0 0 0 0 15 7 0 0 4
432 202
432 121
585 121
585 117
0 4 5 0 0 8320 0 0 11 29 0 4
176 187
176 440
947 440
947 254
3 2 6 0 0 8320 0 6 13 0 0 3
697 138
697 205
780 205
0 2 7 0 0 8320 0 0 6 20 0 4
278 300
278 319
742 319
742 147
2 1 8 0 0 4224 0 5 6 0 0 2
740 129
742 129
0 4 9 0 0 4224 0 0 13 13 0 3
529 355
780 355
780 223
3 4 10 0 0 4224 0 7 14 0 0 3
539 126
539 221
579 221
0 2 11 0 0 4096 0 0 7 19 0 3
512 147
585 147
585 135
1 2 9 0 0 0 0 1 14 0 0 4
495 424
529 424
529 203
579 203
0 4 3 0 0 0 0 0 15 18 0 5
627 195
642 195
642 277
384 277
384 220
3 2 12 0 0 4224 0 10 15 0 0 3
321 96
321 202
384 202
7 1 2 0 0 8320 0 13 10 0 0 3
828 205
828 87
367 87
3 2 13 0 0 8320 0 9 10 0 0 3
467 107
467 105
367 105
7 1 3 0 0 0 0 14 9 0 0 3
627 203
627 98
512 98
2 2 11 0 0 8320 0 8 9 0 0 3
345 300
512 300
512 116
1 1 7 0 0 0 0 2 8 0 0 3
208 297
208 300
309 300
3 3 14 0 0 8320 0 14 13 0 0 3
579 212
579 214
780 214
3 3 14 0 0 0 0 15 14 0 0 3
384 211
384 212
579 212
1 3 14 0 0 0 0 3 15 0 0 3
214 133
214 211
384 211
5 5 5 0 0 0 0 14 13 0 0 3
603 245
603 247
804 247
5 5 5 0 0 0 0 15 14 0 0 3
408 244
408 245
603 245
0 5 5 0 0 0 0 0 15 29 0 3
362 187
362 244
408 244
1 1 5 0 0 0 0 14 13 0 0 3
603 182
603 184
804 184
1 1 5 0 0 0 0 15 14 0 0 3
408 181
408 182
603 182
1 1 5 0 0 0 0 4 15 0 0 4
161 187
367 187
367 181
408 181
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
130 285 173 309
132 287 170 303
5 Input
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
142 121 189 145
146 123 184 139
5 Clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
802 153 819 177
806 154 814 170
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
591 142 610 166
596 144 604 160
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
397 140 414 164
401 142 409 158
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
89 177 127 199
96 180 119 196
3 gnd
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
