CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 86 1918 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 182 457 279
42991634 0
0
6 Title:
5 Name:
0
0
0
80
13 Logic Switch~
5 896 289 0 1 11
0 69
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -13 12 -5
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3175 0 0
2
43435 0
0
13 Logic Switch~
5 139 579 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4411 0 0
2
43435 1
0
13 Logic Switch~
5 138 620 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8285 0 0
2
43435 2
0
13 Logic Switch~
5 139 548 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6178 0 0
2
43435 3
0
13 Logic Switch~
5 140 507 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9911 0 0
2
43435 4
0
13 Logic Switch~
5 483 424 0 10 11
0 73 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7251 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 196 297 0 1 11
0 71
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9851 0 0
2
5.89871e-315 5.26354e-315
0
13 Logic Switch~
5 202 133 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9133 0 0
2
5.89871e-315 5.30499e-315
0
5 4081~
219 428 1829 0 3 22
0 9 10 3
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 22 0
1 U
7576 0 0
2
43435 0
0
8 3-In OR~
219 375 1838 0 4 22
0 12 2 11 10
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U10C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 10 0
1 U
9978 0 0
2
43435 0
0
5 4049~
219 264 1817 0 2 22
0 13 15
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U21C
-14 -19 14 -11
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 21 0
1 U
758 0 0
2
43435 0
0
5 4049~
219 264 1799 0 2 22
0 14 16
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U21B
-14 -19 14 -11
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 21 0
1 U
5351 0 0
2
43435 0
0
5 4081~
219 306 1808 0 3 22
0 16 15 12
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 22 0
1 U
7860 0 0
2
43435 0
0
5 4081~
219 438 1642 0 3 22
0 9 17 4
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 22 0
1 U
8118 0 0
2
43435 0
0
5 4081~
219 460 1410 0 3 22
0 9 18 5
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 22 0
1 U
7363 0 0
2
43435 0
0
5 4071~
219 384 1651 0 3 22
0 20 19 17
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
9572 0 0
2
43435 0
0
5 4049~
219 267 1676 0 2 22
0 11 21
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U21A
-14 -19 14 -11
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 21 0
1 U
3608 0 0
2
43435 0
0
5 4049~
219 268 1667 0 2 22
0 2 22
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19F
-14 -19 14 -11
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 19 0
1 U
8671 0 0
2
43435 0
0
5 4073~
219 310 1676 0 4 22
0 22 21 13 19
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U20A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 20 0
1 U
9832 0 0
2
43435 0
0
5 4049~
219 264 1631 0 2 22
0 11 23
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19E
-14 -19 14 -11
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 19 0
1 U
3630 0 0
2
43435 0
0
5 4049~
219 264 1622 0 2 22
0 2 24
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 19 0
1 U
3159 0 0
2
43435 0
0
5 4073~
219 307 1631 0 4 22
0 24 23 14 20
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 18 0
1 U
7384 0 0
2
43435 0
0
5 4049~
219 171 2019 0 2 22
0 14 77
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 3 19 0
1 U
3933 0 0
2
43435 0
0
5 4049~
219 187 1966 0 2 22
0 13 78
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 2 19 0
1 U
8168 0 0
2
43435 0
0
5 4049~
219 228 1906 0 2 22
0 11 79
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U19A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 1 19 0
1 U
5374 0 0
2
43435 0
0
8 4-In OR~
219 407 1419 0 5 22
0 28 27 26 25 18
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U13B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
7500 0 0
2
5.89871e-315 0
0
5 4073~
219 308 1501 0 4 22
0 2 13 14 25
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 18 0
1 U
4207 0 0
2
5.89871e-315 0
0
5 4073~
219 305 1445 0 4 22
0 11 13 14 26
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 18 0
1 U
3844 0 0
2
5.89871e-315 0
0
5 4049~
219 269 1382 0 2 22
0 13 29
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 17 0
1 U
5174 0 0
2
5.89871e-315 0
0
5 4049~
219 270 1373 0 2 22
0 14 30
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 17 0
1 U
5620 0 0
2
5.89871e-315 0
0
5 4073~
219 312 1382 0 4 22
0 30 29 2 27
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 16 0
1 U
5464 0 0
2
5.89871e-315 0
0
5 4049~
219 266 1340 0 2 22
0 14 31
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 17 0
1 U
5444 0 0
2
5.89871e-315 0
0
5 4049~
219 266 1331 0 2 22
0 13 32
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 17 0
1 U
3975 0 0
2
5.89871e-315 0
0
5 4049~
219 266 1322 0 2 22
0 11 33
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 17 0
1 U
5865 0 0
2
5.89871e-315 0
0
5 4073~
219 309 1331 0 4 22
0 33 32 31 28
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 16 0
1 U
859 0 0
2
5.89871e-315 0
0
5 4081~
219 429 1147 0 3 22
0 9 37 6
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 12 0
1 U
4289 0 0
2
5.89871e-315 0
0
8 3-In OR~
219 375 1156 0 4 22
0 36 35 34 37
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 10 0
1 U
4623 0 0
2
5.89871e-315 0
0
5 4049~
219 262 1214 0 2 22
0 11 38
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 17 0
1 U
9733 0 0
2
5.89871e-315 0
0
5 4049~
219 263 1205 0 2 22
0 2 39
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U14F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 14 0
1 U
4682 0 0
2
5.89871e-315 0
0
5 4073~
219 305 1214 0 4 22
0 39 38 13 34
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 16 0
1 U
8941 0 0
2
5.89871e-315 0
0
5 4049~
219 264 1157 0 2 22
0 2 40
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U14E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 14 0
1 U
3820 0 0
2
5.89871e-315 0
0
5 4049~
219 264 1148 0 2 22
0 13 41
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U14D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 14 0
1 U
8459 0 0
2
5.89871e-315 0
0
5 4073~
219 306 1157 0 4 22
0 41 40 11 35
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 8 0
1 U
3440 0 0
2
5.89871e-315 0
0
5 4070~
219 296 1099 0 3 22
0 13 14 36
0
0 0 624 0
4 4070
-7 -24 21 -16
4 U15A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
5821 0 0
2
5.89871e-315 0
0
5 4081~
219 456 894 0 3 22
0 9 42 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 12 0
1 U
775 0 0
2
5.89871e-315 0
0
8 4-In OR~
219 401 903 0 5 22
0 46 45 44 43 42
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U13A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
8472 0 0
2
5.89871e-315 0
0
5 4049~
219 277 1008 0 2 22
0 14 47
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 11 0
1 U
5642 0 0
2
5.89871e-315 5.30499e-315
0
5 4049~
219 277 990 0 2 22
0 11 48
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 11 0
1 U
5711 0 0
2
5.89871e-315 5.26354e-315
0
5 4081~
219 320 999 0 3 22
0 48 47 43
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
8118 0 0
2
5.89871e-315 0
0
5 4073~
219 319 937 0 4 22
0 11 13 14 44
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 8 0
1 U
3757 0 0
2
5.89871e-315 0
0
5 4081~
219 319 881 0 3 22
0 50 49 45
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U12A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
3882 0 0
2
5.89871e-315 5.30499e-315
0
5 4049~
219 276 872 0 2 22
0 2 50
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 11 0
1 U
9366 0 0
2
5.89871e-315 5.26354e-315
0
5 4049~
219 276 890 0 2 22
0 11 49
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 11 0
1 U
5650 0 0
2
5.89871e-315 0
0
5 4049~
219 276 835 0 2 22
0 13 51
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 11 0
1 U
7718 0 0
2
5.89871e-315 0
0
5 4049~
219 276 817 0 2 22
0 11 52
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 11 0
1 U
6825 0 0
2
5.89871e-315 0
0
5 4081~
219 319 826 0 3 22
0 52 51 46
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
8223 0 0
2
5.89871e-315 0
0
5 4081~
219 576 669 0 3 22
0 9 53 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
4773 0 0
2
5.89871e-315 0
0
8 3-In OR~
219 523 678 0 4 22
0 56 55 54 53
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 10 0
1 U
7329 0 0
2
5.89871e-315 0
0
5 4049~
219 406 737 0 2 22
0 59 60
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 5 0
1 U
5290 0 0
2
43435 6
0
5 4082~
219 449 741 0 5 22
0 2 60 58 57 54
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
6210 0 0
2
43435 7
0
5 4049~
219 420 688 0 2 22
0 57 61
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 5 0
1 U
4522 0 0
2
43435 8
0
5 4073~
219 461 679 0 4 22
0 58 59 61 55
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
4399 0 0
2
43435 9
0
5 4049~
219 421 627 0 2 22
0 58 62
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 5 0
1 U
6836 0 0
2
43435 10
0
5 4081~
219 463 618 0 3 22
0 59 62 56
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
5657 0 0
2
43435 11
0
5 4049~
219 222 226 0 2 22
0 9 64
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 5 0
1 U
3900 0 0
2
5.89871e-315 5.32571e-315
0
5 4081~
219 265 217 0 3 22
0 65 64 63
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
9532 0 0
2
5.89871e-315 5.34643e-315
0
5 4081~
219 236 609 0 3 22
0 9 14 57
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
347 0 0
2
43435 12
0
5 4081~
219 233 569 0 3 22
0 9 13 58
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
8304 0 0
2
43435 13
0
5 4081~
219 234 532 0 3 22
0 9 11 59
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
3414 0 0
2
43435 14
0
5 4049~
219 755 129 0 2 22
0 68 72
0
0 0 624 512
4 4049
-7 -24 21 -16
3 U5B
-5 -20 16 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
4979 0 0
2
5.89871e-315 5.3568e-315
0
5 4081~
219 722 138 0 3 22
0 72 71 70
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4B
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
4312 0 0
2
5.89871e-315 5.36716e-315
0
5 4071~
219 566 126 0 3 22
0 68 2 74
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3B
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
8210 0 0
2
5.89871e-315 5.37752e-315
0
5 4049~
219 324 300 0 2 22
0 71 2
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
8709 0 0
2
5.89871e-315 5.38788e-315
0
5 4081~
219 492 107 0 3 22
0 67 2 76
0
0 0 624 512
4 4081
-7 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
8410 0 0
2
5.89871e-315 5.39306e-315
0
5 4071~
219 348 96 0 3 22
0 66 76 75
0
0 0 624 512
4 4071
-7 -24 21 -16
3 U3A
1 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
6112 0 0
2
5.89871e-315 5.39824e-315
0
12 Hex Display~
7 956 230 0 16 19
10 66 67 68 69 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4562 0 0
2
5.89871e-315 5.40342e-315
0
7 Pulser~
4 150 91 0 10 12
0 80 81 82 83 0 0 5 5 3
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3901 0 0
2
43435 15
0
5 4027~
219 804 241 0 7 32
0 4 70 63 73 3 84 66
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
5761 0 0
2
43435 16
0
5 4027~
219 603 239 0 7 32
0 6 73 63 74 5 85 67
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
510 0 0
2
43435 17
0
5 4027~
219 408 238 0 7 32
0 8 75 63 67 7 86 68
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3190 0 0
2
43435 18
0
146
0 1 2 0 0 4096 0 0 60 2 0 3
350 441
350 728
425 728
0 0 2 0 0 0 0 0 0 145 90 3
350 300
350 442
340 442
3 5 3 0 0 8320 0 9 78 0 0 3
449 1829
804 1829
804 247
3 1 4 0 0 8320 0 14 78 0 0 4
459 1642
848 1642
848 184
804 184
3 5 5 0 0 8320 0 15 79 0 0 4
481 1410
718 1410
718 245
603 245
3 1 6 0 0 8320 0 36 79 0 0 4
450 1147
670 1147
670 182
603 182
3 5 7 0 0 8336 0 45 80 0 0 6
477 894
618 894
618 478
409 478
409 244
408 244
3 1 8 0 0 12416 0 57 80 0 0 5
597 669
597 487
366 487
366 181
408 181
0 1 9 0 0 8192 0 0 9 18 0 4
414 1619
390 1619
390 1820
404 1820
2 4 10 0 0 4224 0 9 10 0 0 2
404 1838
408 1838
0 3 11 0 0 4096 0 0 10 34 0 2
198 1847
362 1847
0 2 2 0 0 8192 0 0 10 26 0 3
40 1667
40 1838
363 1838
3 1 12 0 0 4224 0 13 10 0 0 3
327 1808
362 1808
362 1829
1 0 13 0 0 4096 0 11 0 0 74 2
249 1817
172 1817
1 0 14 0 0 4096 0 12 0 0 75 2
249 1799
157 1799
2 2 15 0 0 4224 0 11 13 0 0 2
285 1817
282 1817
2 1 16 0 0 4224 0 12 13 0 0 2
285 1799
282 1799
0 1 9 0 0 8192 0 0 14 20 0 3
436 1376
414 1376
414 1633
2 3 17 0 0 4224 0 14 16 0 0 2
414 1651
417 1651
0 1 9 0 0 0 0 0 15 59 0 5
405 1089
376 1089
376 1307
436 1307
436 1401
2 5 18 0 0 4224 0 15 26 0 0 2
436 1419
440 1419
4 2 19 0 0 4224 0 19 16 0 0 3
331 1676
371 1676
371 1660
4 1 20 0 0 4224 0 22 16 0 0 3
328 1631
371 1631
371 1642
3 0 13 0 0 4096 0 19 0 0 74 2
286 1685
173 1685
1 0 11 0 0 0 0 17 0 0 73 2
252 1676
198 1676
0 1 2 0 0 0 0 0 18 32 0 3
40 1622
40 1667
253 1667
2 2 21 0 0 4224 0 17 19 0 0 2
288 1676
286 1676
2 1 22 0 0 4224 0 18 19 0 0 2
289 1667
286 1667
3 0 14 0 0 4096 0 22 0 0 75 2
283 1640
157 1640
1 0 11 0 0 0 0 20 0 0 73 2
249 1631
198 1631
2 2 23 0 0 4224 0 20 22 0 0 2
285 1631
283 1631
0 1 2 0 0 0 0 0 21 41 0 3
40 1491
40 1622
249 1622
2 1 24 0 0 4224 0 21 22 0 0 2
285 1622
283 1622
0 1 11 0 0 4096 0 0 25 73 0 3
198 1711
198 1906
213 1906
4 4 25 0 0 8320 0 27 26 0 0 4
329 1501
351 1501
351 1433
390 1433
4 3 26 0 0 8320 0 28 26 0 0 3
326 1445
326 1424
390 1424
4 2 27 0 0 4224 0 31 26 0 0 4
333 1382
379 1382
379 1415
390 1415
4 1 28 0 0 8320 0 35 26 0 0 3
330 1331
390 1331
390 1406
3 0 14 0 0 4096 0 27 0 0 75 2
284 1510
157 1510
2 0 13 0 0 0 0 27 0 0 74 2
284 1501
174 1501
0 1 2 0 0 0 0 0 27 47 0 3
40 1389
40 1492
284 1492
3 0 14 0 0 0 0 28 0 0 75 2
281 1454
157 1454
2 0 13 0 0 0 0 28 0 0 74 2
281 1445
174 1445
1 0 11 0 0 0 0 28 0 0 73 2
281 1436
198 1436
1 0 14 0 0 0 0 30 0 0 75 2
255 1373
158 1373
1 0 13 0 0 0 0 29 0 0 74 2
254 1382
174 1382
0 3 2 0 0 0 0 0 31 63 0 3
40 1204
40 1391
288 1391
2 2 29 0 0 4224 0 29 31 0 0 2
290 1382
288 1382
2 1 30 0 0 4224 0 30 31 0 0 2
291 1373
288 1373
1 0 14 0 0 0 0 32 0 0 75 2
251 1340
158 1340
1 0 13 0 0 0 0 33 0 0 74 2
251 1331
174 1331
0 1 11 0 0 0 0 0 34 73 0 3
199 1321
199 1322
251 1322
2 3 31 0 0 4224 0 32 35 0 0 2
287 1340
285 1340
2 2 32 0 0 4224 0 33 35 0 0 4
287 1331
284 1331
284 1331
285 1331
2 1 33 0 0 4224 0 34 35 0 0 4
287 1322
284 1322
284 1322
285 1322
4 3 34 0 0 4224 0 40 37 0 0 3
326 1214
326 1165
362 1165
4 2 35 0 0 12416 0 43 37 0 0 4
327 1157
336 1157
336 1156
363 1156
3 1 36 0 0 8320 0 44 37 0 0 3
329 1099
362 1099
362 1147
0 1 9 0 0 8192 0 0 36 76 0 3
432 854
405 854
405 1138
2 4 37 0 0 4224 0 36 37 0 0 2
405 1156
408 1156
3 0 13 0 0 0 0 40 0 0 74 2
281 1223
174 1223
1 0 11 0 0 0 0 38 0 0 73 2
247 1214
199 1214
0 1 2 0 0 0 0 0 39 67 0 3
40 1156
40 1205
248 1205
2 2 38 0 0 4224 0 38 40 0 0 2
283 1214
281 1214
2 1 39 0 0 4224 0 39 40 0 0 2
284 1205
281 1205
3 0 11 0 0 0 0 43 0 0 73 2
282 1166
199 1166
0 1 2 0 0 0 0 0 41 90 0 3
40 871
40 1157
249 1157
1 0 13 0 0 0 0 42 0 0 74 2
249 1148
174 1148
2 2 40 0 0 4224 0 41 43 0 0 2
285 1157
282 1157
2 1 41 0 0 4224 0 42 43 0 0 2
285 1148
282 1148
2 0 14 0 0 0 0 44 0 0 75 2
280 1108
158 1108
0 1 13 0 0 0 0 0 44 74 0 3
174 1091
174 1090
280 1090
0 0 11 0 0 16512 0 0 0 86 0 5
196 928
199 928
199 1321
198 1321
198 1716
0 1 13 0 0 4224 0 0 24 87 0 6
174 936
174 1501
173 1501
173 1685
172 1685
172 1966
0 1 14 0 0 12416 0 0 23 88 0 5
158 944
158 1373
157 1373
157 2019
156 2019
0 1 9 0 0 0 0 0 45 97 0 5
552 621
531 621
531 831
432 831
432 885
2 5 42 0 0 4224 0 45 46 0 0 2
432 903
434 903
3 4 43 0 0 8320 0 49 46 0 0 3
341 999
384 999
384 917
4 3 44 0 0 8320 0 50 46 0 0 4
340 937
355 937
355 908
384 908
3 2 45 0 0 4224 0 51 46 0 0 4
340 881
362 881
362 899
384 899
3 1 46 0 0 8320 0 56 46 0 0 3
340 826
384 826
384 890
0 1 14 0 0 0 0 0 47 88 0 3
207 946
207 1008
262 1008
0 1 11 0 0 0 0 0 48 86 0 3
242 928
242 990
262 990
2 2 47 0 0 4224 0 47 49 0 0 2
298 1008
296 1008
2 1 48 0 0 4224 0 48 49 0 0 2
298 990
296 990
0 1 11 0 0 0 0 0 50 94 0 3
196 817
196 928
295 928
0 2 13 0 0 0 0 0 50 93 0 3
174 835
174 937
295 937
0 3 14 0 0 0 0 0 50 126 0 3
158 618
158 946
295 946
0 1 11 0 0 0 0 0 53 94 0 3
231 817
231 890
261 890
0 1 2 0 0 8320 0 0 52 0 0 4
344 442
40 442
40 872
261 872
2 2 49 0 0 4224 0 53 51 0 0 2
297 890
295 890
2 1 50 0 0 4224 0 52 51 0 0 2
297 872
295 872
0 1 13 0 0 0 0 0 54 127 0 3
162 578
162 835
261 835
0 1 11 0 0 0 0 0 55 129 0 3
170 541
170 817
261 817
2 2 51 0 0 4224 0 54 56 0 0 2
297 835
295 835
2 1 52 0 0 4224 0 55 56 0 0 2
297 817
295 817
0 1 9 0 0 4224 0 0 57 130 0 3
203 507
552 507
552 660
2 4 53 0 0 4224 0 57 58 0 0 2
552 678
556 678
5 3 54 0 0 8320 0 60 58 0 0 3
470 741
510 741
510 687
4 2 55 0 0 8320 0 62 58 0 0 3
482 679
482 678
511 678
3 1 56 0 0 8320 0 64 58 0 0 3
484 618
510 618
510 669
0 4 57 0 0 8320 0 0 60 106 0 3
257 688
257 755
425 755
0 3 58 0 0 4096 0 0 60 107 0 3
375 670
375 746
425 746
0 1 59 0 0 8192 0 0 59 105 0 3
332 679
332 737
391 737
0 2 59 0 0 8320 0 0 62 108 0 3
280 532
280 679
437 679
3 1 57 0 0 0 0 67 61 0 0 3
257 609
257 688
405 688
0 1 58 0 0 0 0 0 62 109 0 3
375 627
375 670
437 670
3 1 59 0 0 0 0 69 64 0 0 4
255 532
320 532
320 609
439 609
3 1 58 0 0 12416 0 68 63 0 0 4
254 569
300 569
300 627
406 627
0 1 9 0 0 0 0 0 65 128 0 5
161 507
161 380
84 380
84 226
207 226
2 2 60 0 0 4224 0 59 60 0 0 2
427 737
425 737
2 3 61 0 0 4224 0 61 62 0 0 2
441 688
437 688
2 2 62 0 0 4224 0 63 64 0 0 2
442 627
439 627
3 3 63 0 0 8320 0 79 78 0 0 3
579 212
579 214
780 214
3 3 63 0 0 0 0 80 79 0 0 3
384 211
384 212
579 212
3 3 63 0 0 0 0 66 80 0 0 4
286 217
342 217
342 211
384 211
2 2 64 0 0 4224 0 65 66 0 0 2
243 226
241 226
1 1 65 0 0 8320 0 8 66 0 0 3
214 133
241 133
241 208
0 5 7 0 0 128 0 0 80 0 0 2
408 238
408 244
0 1 66 0 0 12288 0 0 76 124 0 6
1016 391
1016 344
1004 344
1004 272
965 272
965 254
0 2 67 0 0 8320 0 0 76 140 0 8
635 277
635 429
945 429
945 343
936 343
936 319
959 319
959 254
0 3 68 0 0 12416 0 0 76 132 0 9
432 152
456 152
456 470
882 470
882 346
873 346
873 310
953 310
953 254
1 4 69 0 0 8320 0 1 76 0 0 3
908 289
908 254
947 254
0 0 66 0 0 4096 0 0 0 142 0 4
828 139
1085 139
1085 391
1013 391
0 1 9 0 0 0 0 0 67 128 0 3
194 560
194 600
212 600
1 2 14 0 0 0 0 3 67 0 0 3
150 620
150 618
212 618
1 2 13 0 0 0 0 2 68 0 0 3
151 579
151 578
209 578
1 1 9 0 0 0 0 5 68 0 0 4
152 507
176 507
176 560
209 560
1 2 11 0 0 0 0 4 69 0 0 3
151 548
151 541
210 541
0 1 9 0 0 0 0 0 69 128 0 4
174 507
203 507
203 523
210 523
0 1 68 0 0 0 0 0 70 132 0 4
531 121
531 41
776 41
776 129
7 1 68 0 0 0 0 80 72 0 0 4
432 202
432 121
585 121
585 117
3 2 70 0 0 8320 0 71 78 0 0 3
697 138
697 205
780 205
0 2 71 0 0 8320 0 0 71 146 0 4
278 300
278 319
742 319
742 147
2 1 72 0 0 4224 0 70 71 0 0 2
740 129
742 129
0 4 73 0 0 4224 0 0 78 139 0 3
529 355
780 355
780 223
3 4 74 0 0 4224 0 72 79 0 0 3
539 126
539 221
579 221
0 2 2 0 0 0 0 0 72 145 0 3
512 147
585 147
585 135
1 2 73 0 0 0 0 6 79 0 0 4
495 424
529 424
529 203
579 203
0 4 67 0 0 0 0 0 80 144 0 5
627 195
642 195
642 277
384 277
384 220
3 2 75 0 0 4224 0 75 80 0 0 3
321 96
321 202
384 202
7 1 66 0 0 8320 0 78 75 0 0 3
828 205
828 87
367 87
3 2 76 0 0 8320 0 74 75 0 0 3
467 107
467 105
367 105
7 1 67 0 0 0 0 79 74 0 0 3
627 203
627 98
512 98
2 2 2 0 0 128 0 73 74 0 0 3
345 300
512 300
512 116
1 1 71 0 0 0 0 7 73 0 0 3
208 297
208 300
309 300
14
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
122 340 274 364
127 342 268 358
18 1 = multiplos de 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
121 319 273 343
126 321 267 337
18 0 = multiplos de 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
72 539 106 563
77 540 100 556
3 MSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
71 493 125 517
75 495 120 511
6 Ativar
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
397 140 414 164
401 142 409 158
1 X
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
591 142 610 166
596 144 604 160
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
802 153 819 177
806 154 814 170
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
142 121 189 145
146 123 184 139
5 Clock
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
130 285 173 309
132 287 170 303
5 Input
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
484 865 511 889
489 867 505 883
2 R1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
575 629 596 653
577 631 593 647
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
49 851 91 875
54 853 85 869
4 Modo
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
59 1111 133 1135
64 1113 127 1129
8 Q3,Q2,Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
63 1442 137 1466
68 1444 131 1460
8 Q3,Q2,Q1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
