CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 20 1 140 10
176 86 1918 980
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 182 457 279
42991634 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 750 187 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5881 0 0
2
43430.5 0
0
13 Logic Switch~
5 316 392 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3275 0 0
2
43430.5 0
0
13 Logic Switch~
5 863 393 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4203 0 0
2
5.89871e-315 0
0
13 Logic Switch~
5 56 54 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
5.89871e-315 0
0
5 4049~
219 292 581 0 2 22
0 9 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 6 0
1 U
9102 0 0
2
43430.5 0
0
5 4049~
219 226 372 0 2 22
0 4 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 6 0
1 U
5586 0 0
2
43430.5 0
0
5 4049~
219 213 349 0 2 22
0 4 12
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 6 0
1 U
525 0 0
2
43430.5 0
0
5 4049~
219 214 331 0 2 22
0 9 13
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U6B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 6 0
1 U
6206 0 0
2
43430.5 0
0
5 4081~
219 257 340 0 3 22
0 13 12 11
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3418 0 0
2
43430.5 0
0
5 4081~
219 190 221 0 3 22
0 5 3 14
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
9312 0 0
2
43430.5 0
0
9 CC 7-Seg~
183 781 258 0 17 19
10 5 4 4 3 6 6 5 16 2
0 0 0 0 1 1 0 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
7419 0 0
2
5.89871e-315 0
0
5 4027~
219 420 482 0 7 32
0 15 3 7 3 15 26 4
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
472 0 0
2
5.89871e-315 5.26354e-315
0
5 4027~
219 419 599 0 7 32
0 15 5 7 8 15 27 3
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
4714 0 0
2
5.89871e-315 0
0
5 4027~
219 418 368 0 7 32
0 15 11 7 10 15 28 5
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
9386 0 0
2
5.89871e-315 0
0
5 4027~
219 419 251 0 7 32
0 15 14 7 3 15 29 9
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
7610 0 0
2
5.89871e-315 0
0
36
1 9 2 0 0 8320 0 1 11 0 0 3
762 187
781 187
781 216
0 4 3 0 0 8192 0 0 11 27 0 3
579 569
778 569
778 294
0 3 4 0 0 8192 0 0 11 4 0 3
765 446
772 446
772 294
0 2 4 0 0 0 0 0 11 21 0 3
620 446
766 446
766 294
0 7 5 0 0 8192 0 0 11 6 0 3
760 332
796 332
796 294
0 1 5 0 0 4096 0 0 11 28 0 3
580 332
760 332
760 294
0 5 6 0 0 8192 0 0 11 8 0 3
790 353
784 353
784 294
1 6 6 0 0 8320 0 3 11 0 0 4
875 393
875 353
790 353
790 294
0 3 7 0 0 8192 0 0 13 10 0 3
68 455
68 572
395 572
0 3 7 0 0 8320 0 0 12 11 0 3
68 339
68 455
396 455
0 3 7 0 0 0 0 0 14 12 0 3
68 224
68 341
394 341
1 3 7 0 0 0 0 4 15 0 0 3
68 54
68 224
395 224
2 4 8 0 0 4224 0 5 13 0 0 2
313 581
395 581
0 1 9 0 0 4096 0 0 5 22 0 3
141 331
141 581
277 581
0 2 5 0 0 8192 0 0 13 28 0 5
544 332
544 514
276 514
276 563
395 563
4 0 3 0 0 0 0 12 0 0 27 2
396 464
166 464
2 0 3 0 0 0 0 12 0 0 27 2
396 446
166 446
2 4 10 0 0 12416 0 6 14 0 0 4
247 372
287 372
287 350
394 350
1 0 4 0 0 0 0 6 0 0 21 2
211 372
116 372
3 2 11 0 0 8320 0 9 14 0 0 3
278 340
278 332
394 332
7 1 4 0 0 12416 0 12 7 0 0 6
444 446
622 446
622 641
116 641
116 349
198 349
7 1 9 0 0 8320 0 15 8 0 0 5
443 215
443 60
116 60
116 331
199 331
2 2 12 0 0 4224 0 7 9 0 0 2
234 349
233 349
2 1 13 0 0 4224 0 8 9 0 0 2
235 331
233 331
0 4 3 0 0 0 0 0 15 27 0 4
166 249
222 249
222 233
395 233
3 2 14 0 0 12416 0 10 15 0 0 4
211 221
219 221
219 215
395 215
7 2 3 0 0 12416 0 13 10 0 0 5
443 563
579 563
579 631
166 631
166 230
7 1 5 0 0 12416 0 14 10 0 0 5
442 332
580 332
580 101
166 101
166 212
0 5 15 0 0 8192 0 0 13 30 0 3
328 541
328 605
419 605
0 1 15 0 0 0 0 0 13 31 0 3
328 488
328 542
419 542
0 5 15 0 0 8192 0 0 12 32 0 3
328 423
328 488
420 488
1 1 15 0 0 0 0 2 12 0 0 3
328 392
328 425
420 425
0 5 15 0 0 0 0 0 14 36 0 3
328 371
328 374
418 374
0 1 15 0 0 0 0 0 14 36 0 3
328 312
328 311
418 311
0 5 15 0 0 0 0 0 15 36 0 3
328 254
328 257
419 257
1 1 15 0 0 4224 0 2 15 0 0 3
328 392
328 194
419 194
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
494 539 513 563
499 541 507 557
1 W
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
485 430 504 454
490 432 498 448
1 Z
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
484 318 503 342
489 320 497 336
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
484 175 503 199
489 177 497 193
1 X
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
