CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 140 10
176 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
47
13 Logic Switch~
5 106 95 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 I
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43402.8 0
0
13 Logic Switch~
5 278 88 0 1 11
0 2
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89865e-315 0
0
13 Logic Switch~
5 241 94 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89865e-315 0
0
13 Logic Switch~
5 192 92 0 1 11
0 20
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89865e-315 5.26354e-315
0
13 Logic Switch~
5 148 93 0 1 11
0 36
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89865e-315 5.30499e-315
0
8 2-In OR~
219 496 946 0 3 22
0 4 3 43
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 33 0
1 U
5572 0 0
2
43402.9 0
0
9 2-In AND~
219 461 987 0 3 22
0 5 6 3
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 34 0
1 U
8901 0 0
2
43402.9 0
0
5 4030~
219 402 974 0 3 22
0 7 7 5
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 35 0
1 U
7361 0 0
2
43402.9 0
0
9 2-In AND~
219 385 913 0 3 22
0 8 7 4
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 34 0
1 U
4747 0 0
2
43402.9 0
0
5 4049~
219 334 902 0 2 22
0 6 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 29 0
1 U
972 0 0
2
43402.9 0
0
8 2-In OR~
219 740 748 0 3 22
0 10 9 44
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 33 0
1 U
3472 0 0
2
43402.9 0
0
9 2-In AND~
219 684 839 0 3 22
0 11 6 9
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 34 0
1 U
9998 0 0
2
43402.9 0
0
8 2-In OR~
219 611 799 0 3 22
0 13 12 11
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
3536 0 0
2
43402.9 0
0
8 2-In OR~
219 514 761 0 3 22
0 15 14 13
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U8A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
4597 0 0
2
43402.9 0
0
9 2-In AND~
219 453 729 0 3 22
0 20 16 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
3835 0 0
2
43402.9 0
0
9 2-In AND~
219 381 732 0 3 22
0 18 17 16
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
3670 0 0
2
43402.9 0
0
9 2-In AND~
219 448 789 0 3 22
0 19 7 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
5616 0 0
2
43402.9 0
0
9 2-In AND~
219 448 839 0 3 22
0 19 2 12
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
9323 0 0
2
43402.9 0
0
5 4049~
219 329 781 0 2 22
0 20 19
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 29 0
1 U
317 0 0
2
43402.9 0
0
5 4049~
219 329 741 0 2 22
0 2 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 29 0
1 U
3108 0 0
2
43402.9 0
0
5 4049~
219 329 722 0 2 22
0 7 18
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 29 0
1 U
4299 0 0
2
43402.9 0
0
9 2-In AND~
219 380 646 0 3 22
0 21 20 10
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
9672 0 0
2
43402.9 0
0
5 4049~
219 323 634 0 2 22
0 6 21
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 29 0
1 U
7876 0 0
2
43402.9 0
0
8 2-In OR~
219 923 421 0 3 22
0 23 22 45
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 31 0
1 U
6369 0 0
2
43402.8 0
0
9 2-In AND~
219 866 526 0 3 22
0 24 6 22
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
9172 0 0
2
43402.8 0
0
8 2-In OR~
219 761 466 0 3 22
0 26 25 24
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
7100 0 0
2
43402.8 0
0
8 2-In OR~
219 649 498 0 3 22
0 28 27 25
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
3820 0 0
2
43402.8 0
0
8 2-In OR~
219 649 391 0 3 22
0 30 29 26
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U6A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
7678 0 0
2
43402.8 0
0
9 2-In AND~
219 592 541 0 3 22
0 32 31 27
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
961 0 0
2
43402.8 0
0
9 2-In AND~
219 540 575 0 3 22
0 33 36 31
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
3178 0 0
2
43402.8 0
0
9 2-In AND~
219 538 522 0 3 22
0 34 35 32
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
3409 0 0
2
43402.8 0
0
5 4049~
219 479 562 0 2 22
0 2 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 29 0
1 U
3951 0 0
2
43402.8 0
0
5 4049~
219 481 534 0 2 22
0 7 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 23 0
1 U
8885 0 0
2
43402.8 0
0
5 4049~
219 479 511 0 2 22
0 20 34
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 23 0
1 U
3780 0 0
2
43402.8 0
0
9 2-In AND~
219 483 463 0 3 22
0 37 2 28
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
9265 0 0
2
43402.8 0
0
9 2-In AND~
219 484 415 0 3 22
0 37 7 29
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
9442 0 0
2
43402.8 0
0
9 2-In AND~
219 485 358 0 3 22
0 37 20 30
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
9424 0 0
2
43402.8 0
0
5 4049~
219 352 344 0 2 22
0 36 37
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 23 0
1 U
9968 0 0
2
43402.8 0
0
9 2-In AND~
219 404 289 0 3 22
0 38 36 23
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
9281 0 0
2
43402.8 0
0
5 4049~
219 352 271 0 2 22
0 6 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 23 0
1 U
8464 0 0
2
43402.8 0
0
9 2-In AND~
219 562 135 0 3 22
0 6 40 39
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
7168 0 0
2
43402.8 0
0
8 2-In OR~
219 482 185 0 3 22
0 42 41 40
0
0 0 624 0
5 74F32
-18 -24 17 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
3171 0 0
2
43402.8 0
0
8 2-In OR~
219 400 205 0 3 22
0 7 2 41
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U18D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
4139 0 0
2
43402.8 0
0
8 2-In OR~
219 401 168 0 3 22
0 36 20 42
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U18C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
6435 0 0
2
43402.8 0
0
8 2-In OR~
219 1083 719 0 3 22
0 46 47 48
0
0 0 624 0
5 74F32
-18 -24 17 -16
4 U18B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 27 0
1 U
5283 0 0
2
5.89865e-315 5.32571e-315
0
9 2-In AND~
219 1090 769 0 3 22
0 49 50 51
0
0 0 624 0
5 74F08
-18 -24 17 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 26 0
1 U
6874 0 0
2
5.89865e-315 5.34643e-315
0
5 4049~
219 1093 674 0 2 22
0 52 53
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 512 6 2 23 0
1 U
5305 0 0
2
5.89865e-315 5.3568e-315
0
75
0 0 2 0 0 4096 0 0 0 73 0 2
277 1036
526 1036
2 3 3 0 0 8320 0 6 7 0 0 3
483 955
482 955
482 987
1 3 4 0 0 8320 0 6 9 0 0 3
483 937
483 913
406 913
1 3 5 0 0 4224 0 7 8 0 0 3
437 978
437 974
435 974
0 2 6 0 0 4096 0 0 7 71 0 3
106 1002
437 1002
437 996
2 0 7 0 0 4096 0 8 0 0 74 2
386 983
241 983
1 0 7 0 0 0 0 8 0 0 74 2
386 965
241 965
1 2 8 0 0 8320 0 9 10 0 0 3
361 904
361 902
355 902
0 2 7 0 0 0 0 0 9 74 0 3
241 925
361 925
361 922
0 1 6 0 0 0 0 0 10 71 0 3
106 903
319 903
319 902
2 3 9 0 0 4224 0 11 12 0 0 3
727 757
727 839
705 839
1 3 10 0 0 8320 0 11 22 0 0 3
727 739
727 646
401 646
1 3 11 0 0 4224 0 12 13 0 0 4
660 830
660 814
644 814
644 799
0 2 6 0 0 4096 0 0 12 71 0 3
106 872
660 872
660 848
2 3 12 0 0 4224 0 13 18 0 0 3
598 808
469 808
469 839
1 3 13 0 0 8320 0 13 14 0 0 3
598 790
598 761
547 761
2 3 14 0 0 8320 0 14 17 0 0 3
501 770
501 789
469 789
1 3 15 0 0 4224 0 14 15 0 0 3
501 752
474 752
474 729
3 2 16 0 0 8320 0 16 15 0 0 3
402 732
402 738
429 738
2 2 17 0 0 4224 0 16 20 0 0 2
357 741
350 741
1 2 18 0 0 8320 0 16 21 0 0 3
357 723
357 722
350 722
0 2 2 0 0 0 0 0 18 73 0 3
277 851
424 851
424 848
0 1 19 0 0 8192 0 0 18 24 0 3
366 781
366 830
424 830
2 1 19 0 0 4224 0 19 17 0 0 3
350 781
424 781
424 780
0 2 7 0 0 4096 0 0 17 74 0 3
241 801
424 801
424 798
0 1 20 0 0 4096 0 0 19 72 0 2
192 781
314 781
0 1 2 0 0 0 0 0 20 73 0 2
277 741
314 741
0 1 7 0 0 0 0 0 21 74 0 2
241 722
314 722
0 1 20 0 0 4096 0 0 15 72 0 3
192 706
429 706
429 720
1 2 21 0 0 4224 0 22 23 0 0 3
356 637
344 637
344 634
0 2 20 0 0 0 0 0 22 72 0 4
192 659
207 659
207 655
356 655
0 1 6 0 0 0 0 0 23 71 0 2
106 634
308 634
2 3 22 0 0 8320 0 24 25 0 0 3
910 430
887 430
887 526
1 3 23 0 0 8320 0 24 39 0 0 3
910 412
910 289
425 289
1 3 24 0 0 4224 0 25 26 0 0 3
842 517
842 466
794 466
0 2 6 0 0 4096 0 0 25 71 0 3
106 614
842 614
842 535
2 3 25 0 0 8320 0 26 27 0 0 3
748 475
748 498
682 498
1 3 26 0 0 4224 0 26 28 0 0 3
748 457
682 457
682 391
2 3 27 0 0 8320 0 27 29 0 0 3
636 507
613 507
613 541
1 3 28 0 0 4224 0 27 35 0 0 4
636 489
519 489
519 463
504 463
2 3 29 0 0 4224 0 28 36 0 0 3
636 400
505 400
505 415
1 3 30 0 0 8320 0 28 37 0 0 4
636 382
636 373
506 373
506 358
2 3 31 0 0 4224 0 29 30 0 0 3
568 550
568 575
561 575
3 1 32 0 0 4224 0 31 29 0 0 3
559 522
559 532
568 532
1 2 33 0 0 8320 0 30 32 0 0 3
516 566
516 562
500 562
1 2 34 0 0 8320 0 31 34 0 0 3
514 513
514 511
500 511
2 2 35 0 0 4224 0 31 33 0 0 3
514 531
502 531
502 534
0 2 36 0 0 4096 0 0 30 75 0 3
148 588
516 588
516 584
0 1 2 0 0 0 0 0 32 73 0 2
277 562
464 562
0 1 7 0 0 4096 0 0 33 74 0 2
241 534
466 534
0 1 20 0 0 4096 0 0 34 72 0 2
192 511
464 511
0 2 2 0 0 0 0 0 35 73 0 2
277 472
459 472
0 1 37 0 0 4224 0 0 35 56 0 3
413 344
413 454
459 454
0 2 7 0 0 0 0 0 36 74 0 3
241 426
460 426
460 424
0 1 37 0 0 0 0 0 36 56 0 4
386 344
386 405
460 405
460 406
2 1 37 0 0 0 0 38 37 0 0 3
373 344
461 344
461 349
0 2 20 0 0 0 0 0 37 72 0 3
192 372
461 372
461 367
0 1 36 0 0 0 0 0 38 75 0 2
148 344
337 344
2 0 36 0 0 0 0 39 0 0 75 2
380 298
148 298
1 2 38 0 0 4224 0 39 40 0 0 3
380 280
380 271
373 271
0 1 6 0 0 0 0 0 40 71 0 2
106 271
337 271
3 0 39 0 0 4224 0 41 0 0 0 2
583 135
618 135
1 0 6 0 0 0 0 41 0 0 71 2
538 126
106 126
2 3 40 0 0 8320 0 41 42 0 0 3
538 144
515 144
515 185
2 3 41 0 0 8320 0 42 43 0 0 3
469 194
469 205
433 205
1 3 42 0 0 8320 0 42 44 0 0 3
469 176
469 168
434 168
2 0 2 0 0 0 0 43 0 0 73 2
387 214
277 214
1 0 7 0 0 0 0 43 0 0 74 2
387 196
241 196
2 0 20 0 0 0 0 44 0 0 72 2
388 177
192 177
1 0 36 0 0 0 0 44 0 0 75 2
388 159
148 159
1 0 6 0 0 4224 0 1 0 0 0 3
106 107
106 2172
125 2172
0 1 20 0 0 8320 0 0 4 0 0 3
190 2189
192 2189
192 104
1 0 2 0 0 8320 0 2 0 0 0 4
278 100
277 100
277 2179
300 2179
1 0 7 0 0 4224 0 3 0 0 0 3
241 106
241 2185
264 2185
1 0 36 0 0 4224 0 5 0 0 0 3
148 105
148 2187
166 2187
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
536 1029 558 1053
543 1034 550 1050
1 J
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
530 930 552 954
537 936 544 952
1 H
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
780 738 802 762
787 743 794 759
1 G
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
954 401 976 425
961 407 968 423
1 F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
618 121 640 145
625 126 632 142
1 E
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
