CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1918 996
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
5 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 925 163 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3907 0 0
2
43402.7 4
0
13 Logic Switch~
5 817 163 0 1 11
0 28
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4389 0 0
2
43402.7 3
0
13 Logic Switch~
5 724 152 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7762 0 0
2
43402.7 2
0
13 Logic Switch~
5 620 152 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6723 0 0
2
43402.7 1
0
13 Logic Switch~
5 552 149 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6871 0 0
2
43402.7 0
0
13 Logic Switch~
5 46 145 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4198 0 0
2
43402.7 4
0
13 Logic Switch~
5 135 144 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
970 0 0
2
43402.7 3
0
13 Logic Switch~
5 239 144 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
319 0 0
2
43402.7 2
0
13 Logic Switch~
5 332 155 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3663 0 0
2
43402.7 1
0
13 Logic Switch~
5 440 155 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3512 0 0
2
43402.7 0
0
14 Logic Display~
6 1742 872 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7555 0 0
2
43402.8 0
0
14 Logic Display~
6 1736 805 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9776 0 0
2
43402.8 0
0
14 Logic Display~
6 1729 727 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6596 0 0
2
43402.8 0
0
14 Logic Display~
6 1728 661 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6750 0 0
2
43402.8 0
0
14 Logic Display~
6 1907 1109 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9636 0 0
2
43402.8 0
0
5 4069~
219 1565 1156 0 2 22
0 10 9
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U6A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
5369 0 0
2
43402.8 0
0
6 74LS83
105 1775 1111 0 14 29
0 2 2 2 12 2 2 2 11 9
30 31 32 8 33
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U5
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 0 0 0 0
1 U
8555 0 0
2
43402.7 0
0
5 4081~
219 1686 896 0 3 22
0 16 10 7
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
4690 0 0
2
43402.7 0
0
5 4081~
219 1682 821 0 3 22
0 15 10 6
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
9145 0 0
2
43402.7 0
0
5 4081~
219 1681 742 0 3 22
0 14 10 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
5246 0 0
2
43402.7 0
0
5 4081~
219 1676 679 0 3 22
0 13 10 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9111 0 0
2
43402.7 0
0
7 Ground~
168 1224 853 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6717 0 0
2
43402.7 0
0
6 74LS83
105 1505 782 0 14 29
0 23 22 21 3 17 18 19 20 2
13 14 15 16 10
0
0 0 4848 0
5 74F83
-18 -60 17 -52
2 U3
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 0 0 0 0
1 U
3487 0 0
2
43402.7 0
0
5 4030~
219 1143 402 0 3 22
0 3 28 21
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9604 0 0
2
43402.7 15
0
5 4030~
219 1276 501 0 3 22
0 24 27 22
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3921 0 0
2
43402.7 14
0
5 4030~
219 1403 607 0 3 22
0 26 25 23
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
8146 0 0
2
43402.7 13
0
5 4071~
219 1073 485 0 3 22
0 28 3 24
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4506 0 0
2
43402.7 11
0
5 4071~
219 1164 576 0 3 22
0 27 24 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U2C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
5386 0 0
2
43402.7 10
0
14 Logic Display~
6 1097 263 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7847 0 0
2
43402.7 8
0
14 Logic Display~
6 1213 376 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9261 0 0
2
43402.7 7
0
14 Logic Display~
6 1357 476 0 1 2
10 22
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8231 0 0
2
43402.7 6
0
14 Logic Display~
6 1472 592 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3756 0 0
2
43402.7 5
0
54
0 0 3 0 0 8192 0 0 0 51 40 3
974 304
974 303
1035 303
0 1 2 0 0 4096 0 0 22 27 0 3
1280 835
1224 835
1224 847
3 1 4 0 0 4224 0 21 14 0 0 2
1697 679
1728 679
3 1 5 0 0 8320 0 20 13 0 0 3
1702 742
1702 745
1729 745
3 1 6 0 0 8320 0 19 12 0 0 3
1703 821
1703 823
1736 823
3 1 7 0 0 4224 0 18 11 0 0 3
1707 896
1742 896
1742 890
13 1 8 0 0 8320 0 17 15 0 0 3
1807 1129
1807 1127
1907 1127
2 9 9 0 0 4224 0 16 17 0 0 2
1586 1156
1743 1156
0 1 10 0 0 4224 0 0 16 26 0 3
1544 827
1544 1156
1550 1156
0 8 11 0 0 8320 0 0 17 11 0 3
560 284
560 1138
1743 1138
1 0 11 0 0 0 0 5 0 0 0 3
564 149
560 149
560 299
1 4 12 0 0 8320 0 6 17 0 0 3
58 145
58 1102
1743 1102
0 7 2 0 0 8320 0 0 17 14 0 3
1454 1120
1454 1129
1743 1129
0 6 2 0 0 0 0 0 17 15 0 3
1454 1111
1454 1120
1743 1120
0 5 2 0 0 0 0 0 17 16 0 3
1454 1093
1454 1111
1743 1111
0 3 2 0 0 0 0 0 17 17 0 3
1454 1083
1454 1093
1743 1093
0 2 2 0 0 0 0 0 17 18 0 3
1454 1075
1454 1084
1743 1084
0 1 2 0 0 0 0 0 17 27 0 3
1454 835
1454 1075
1743 1075
10 1 13 0 0 8320 0 23 21 0 0 4
1537 773
1594 773
1594 670
1652 670
0 2 10 0 0 0 0 0 21 22 0 3
1626 751
1626 688
1652 688
11 1 14 0 0 4224 0 23 20 0 0 4
1537 782
1608 782
1608 733
1657 733
0 2 10 0 0 0 0 0 20 24 0 3
1620 830
1620 751
1657 751
12 1 15 0 0 4224 0 23 19 0 0 4
1537 791
1632 791
1632 812
1658 812
0 2 10 0 0 0 0 0 19 26 0 3
1573 827
1573 830
1658 830
13 1 16 0 0 8320 0 23 18 0 0 4
1537 800
1580 800
1580 887
1662 887
14 2 10 0 0 0 0 23 18 0 0 4
1537 827
1573 827
1573 905
1662 905
0 9 2 0 0 0 0 0 23 0 0 3
1264 835
1473 835
1473 827
1 5 17 0 0 8320 0 7 23 0 0 3
147 144
147 782
1473 782
1 6 18 0 0 8320 0 8 23 0 0 3
251 144
251 791
1473 791
1 7 19 0 0 8320 0 9 23 0 0 3
344 155
344 800
1473 800
1 8 20 0 0 8320 0 10 23 0 0 3
452 155
452 809
1473 809
0 4 3 0 0 4224 0 0 23 40 0 3
1060 303
1060 773
1473 773
0 3 21 0 0 4224 0 0 23 39 0 3
1186 402
1186 764
1473 764
0 2 22 0 0 4224 0 0 23 38 0 3
1331 501
1331 755
1473 755
0 1 23 0 0 4224 0 0 23 37 0 3
1441 610
1441 746
1473 746
0 3 24 0 0 4096 0 0 27 46 0 2
1113 485
1106 485
3 1 23 0 0 0 0 26 32 0 0 3
1436 607
1436 610
1472 610
3 1 22 0 0 0 0 25 31 0 0 3
1309 501
1357 501
1357 494
3 1 21 0 0 0 0 24 30 0 0 3
1176 402
1213 402
1213 394
0 1 3 0 0 0 0 0 29 0 0 3
1032 303
1097 303
1097 281
1 2 25 0 0 8320 0 4 26 0 0 3
632 152
632 616
1387 616
3 1 26 0 0 4224 0 28 26 0 0 4
1197 576
1323 576
1323 598
1387 598
0 2 24 0 0 4096 0 0 28 46 0 3
1117 485
1117 585
1151 585
0 1 27 0 0 8192 0 0 28 45 0 3
1023 510
1023 567
1151 567
1 2 27 0 0 8320 0 3 25 0 0 3
736 152
736 510
1260 510
0 1 24 0 0 4224 0 0 25 0 0 4
1109 485
1254 485
1254 492
1260 492
0 2 3 0 0 128 0 0 27 50 0 3
1048 393
1048 494
1060 494
0 1 28 0 0 8192 0 0 27 49 0 3
829 410
829 476
1060 476
1 2 28 0 0 8320 0 2 24 0 0 3
829 163
829 411
1127 411
0 1 3 0 0 0 0 0 24 0 0 3
1043 390
1043 393
1127 393
1 0 3 0 0 0 0 1 0 0 47 5
937 163
974 163
974 381
1048 381
1048 393
0 1 25 0 0 0 0 0 4 0 0 3
635 164
635 152
632 152
0 1 17 0 0 0 0 0 7 0 0 3
150 156
150 144
147 144
0 0 29 0 0 4224 0 0 0 0 0 2
128 1155
128 1138
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
72 58 150 79
77 61 144 76
9 questao 2
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
